module position_cache_to_PE_mapping
#(
	parameter NUM_CELLS = 64, 
	parameter OFFSET_WIDTH = 29, 
	parameter POS_CACHE_WIDTH = 3*OFFSET_WIDTH, 
	parameter NUM_NEIGHBOR_CELLS = 13
)
(
	input [NUM_CELLS*POS_CACHE_WIDTH-1:0] rd_nb_position, 
	input [NUM_CELLS-1:0] broadcast_done, 
	
	output [(NUM_NEIGHBOR_CELLS+1)*NUM_CELLS*POS_CACHE_WIDTH-1:0] rd_nb_position_splitted, 
	output [(NUM_NEIGHBOR_CELLS+1)*NUM_CELLS-1:0] broadcast_done_splitted
);

assign rd_nb_position_splitted[(0*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(0*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[1*POS_CACHE_WIDTH-1:0*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(0*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(0*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[50*POS_CACHE_WIDTH-1:49*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(0*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(0*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[21*POS_CACHE_WIDTH-1:20*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(0*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(0*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[16*POS_CACHE_WIDTH-1:15*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(0*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(0*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[56*POS_CACHE_WIDTH-1:55*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(0*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(0*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[24*POS_CACHE_WIDTH-1:23*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(0*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(0*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[32*POS_CACHE_WIDTH-1:31*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(0*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(0*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[64*POS_CACHE_WIDTH-1:63*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(0*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(0*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[52*POS_CACHE_WIDTH-1:51*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(0*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(0*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[8*POS_CACHE_WIDTH-1:7*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(0*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(0*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[53*POS_CACHE_WIDTH-1:52*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(0*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(0*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[17*POS_CACHE_WIDTH-1:16*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(0*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(0*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[13*POS_CACHE_WIDTH-1:12*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(0*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(0*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[2*POS_CACHE_WIDTH-1:1*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(1*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(1*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[2*POS_CACHE_WIDTH-1:1*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(1*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(1*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[51*POS_CACHE_WIDTH-1:50*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(1*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(1*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[22*POS_CACHE_WIDTH-1:21*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(1*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(1*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[13*POS_CACHE_WIDTH-1:12*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(1*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(1*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[53*POS_CACHE_WIDTH-1:52*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(1*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(1*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[21*POS_CACHE_WIDTH-1:20*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(1*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(1*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[29*POS_CACHE_WIDTH-1:28*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(1*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(1*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[61*POS_CACHE_WIDTH-1:60*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(1*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(1*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[49*POS_CACHE_WIDTH-1:48*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(1*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(1*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[5*POS_CACHE_WIDTH-1:4*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(1*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(1*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[54*POS_CACHE_WIDTH-1:53*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(1*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(1*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[18*POS_CACHE_WIDTH-1:17*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(1*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(1*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[14*POS_CACHE_WIDTH-1:13*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(1*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(1*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[3*POS_CACHE_WIDTH-1:2*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(2*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(2*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[3*POS_CACHE_WIDTH-1:2*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(2*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(2*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[52*POS_CACHE_WIDTH-1:51*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(2*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(2*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[23*POS_CACHE_WIDTH-1:22*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(2*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(2*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[14*POS_CACHE_WIDTH-1:13*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(2*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(2*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[54*POS_CACHE_WIDTH-1:53*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(2*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(2*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[22*POS_CACHE_WIDTH-1:21*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(2*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(2*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[30*POS_CACHE_WIDTH-1:29*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(2*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(2*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[62*POS_CACHE_WIDTH-1:61*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(2*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(2*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[50*POS_CACHE_WIDTH-1:49*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(2*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(2*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[6*POS_CACHE_WIDTH-1:5*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(2*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(2*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[55*POS_CACHE_WIDTH-1:54*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(2*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(2*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[19*POS_CACHE_WIDTH-1:18*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(2*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(2*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[15*POS_CACHE_WIDTH-1:14*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(2*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(2*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[4*POS_CACHE_WIDTH-1:3*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(3*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(3*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[4*POS_CACHE_WIDTH-1:3*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(3*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(3*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[49*POS_CACHE_WIDTH-1:48*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(3*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(3*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[24*POS_CACHE_WIDTH-1:23*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(3*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(3*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[15*POS_CACHE_WIDTH-1:14*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(3*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(3*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[55*POS_CACHE_WIDTH-1:54*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(3*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(3*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[23*POS_CACHE_WIDTH-1:22*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(3*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(3*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[31*POS_CACHE_WIDTH-1:30*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(3*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(3*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[63*POS_CACHE_WIDTH-1:62*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(3*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(3*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[51*POS_CACHE_WIDTH-1:50*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(3*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(3*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[7*POS_CACHE_WIDTH-1:6*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(3*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(3*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[56*POS_CACHE_WIDTH-1:55*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(3*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(3*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[20*POS_CACHE_WIDTH-1:19*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(3*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(3*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[16*POS_CACHE_WIDTH-1:15*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(3*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(3*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[1*POS_CACHE_WIDTH-1:0*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(4*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(4*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[5*POS_CACHE_WIDTH-1:4*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(4*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(4*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[54*POS_CACHE_WIDTH-1:53*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(4*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(4*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[25*POS_CACHE_WIDTH-1:24*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(4*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(4*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[4*POS_CACHE_WIDTH-1:3*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(4*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(4*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[60*POS_CACHE_WIDTH-1:59*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(4*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(4*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[28*POS_CACHE_WIDTH-1:27*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(4*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(4*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[20*POS_CACHE_WIDTH-1:19*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(4*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(4*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[52*POS_CACHE_WIDTH-1:51*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(4*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(4*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[56*POS_CACHE_WIDTH-1:55*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(4*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(4*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[12*POS_CACHE_WIDTH-1:11*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(4*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(4*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[57*POS_CACHE_WIDTH-1:56*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(4*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(4*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[21*POS_CACHE_WIDTH-1:20*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(4*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(4*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[1*POS_CACHE_WIDTH-1:0*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(4*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(4*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[6*POS_CACHE_WIDTH-1:5*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(5*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(5*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[6*POS_CACHE_WIDTH-1:5*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(5*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(5*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[55*POS_CACHE_WIDTH-1:54*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(5*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(5*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[26*POS_CACHE_WIDTH-1:25*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(5*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(5*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[1*POS_CACHE_WIDTH-1:0*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(5*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(5*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[57*POS_CACHE_WIDTH-1:56*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(5*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(5*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[25*POS_CACHE_WIDTH-1:24*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(5*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(5*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[17*POS_CACHE_WIDTH-1:16*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(5*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(5*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[49*POS_CACHE_WIDTH-1:48*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(5*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(5*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[53*POS_CACHE_WIDTH-1:52*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(5*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(5*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[9*POS_CACHE_WIDTH-1:8*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(5*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(5*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[58*POS_CACHE_WIDTH-1:57*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(5*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(5*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[22*POS_CACHE_WIDTH-1:21*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(5*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(5*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[2*POS_CACHE_WIDTH-1:1*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(5*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(5*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[7*POS_CACHE_WIDTH-1:6*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(6*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(6*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[7*POS_CACHE_WIDTH-1:6*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(6*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(6*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[56*POS_CACHE_WIDTH-1:55*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(6*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(6*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[27*POS_CACHE_WIDTH-1:26*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(6*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(6*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[2*POS_CACHE_WIDTH-1:1*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(6*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(6*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[58*POS_CACHE_WIDTH-1:57*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(6*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(6*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[26*POS_CACHE_WIDTH-1:25*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(6*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(6*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[18*POS_CACHE_WIDTH-1:17*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(6*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(6*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[50*POS_CACHE_WIDTH-1:49*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(6*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(6*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[54*POS_CACHE_WIDTH-1:53*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(6*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(6*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[10*POS_CACHE_WIDTH-1:9*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(6*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(6*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[59*POS_CACHE_WIDTH-1:58*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(6*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(6*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[23*POS_CACHE_WIDTH-1:22*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(6*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(6*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[3*POS_CACHE_WIDTH-1:2*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(6*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(6*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[8*POS_CACHE_WIDTH-1:7*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(7*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(7*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[8*POS_CACHE_WIDTH-1:7*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(7*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(7*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[53*POS_CACHE_WIDTH-1:52*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(7*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(7*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[28*POS_CACHE_WIDTH-1:27*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(7*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(7*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[3*POS_CACHE_WIDTH-1:2*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(7*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(7*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[59*POS_CACHE_WIDTH-1:58*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(7*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(7*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[27*POS_CACHE_WIDTH-1:26*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(7*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(7*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[19*POS_CACHE_WIDTH-1:18*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(7*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(7*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[51*POS_CACHE_WIDTH-1:50*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(7*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(7*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[55*POS_CACHE_WIDTH-1:54*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(7*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(7*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[11*POS_CACHE_WIDTH-1:10*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(7*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(7*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[60*POS_CACHE_WIDTH-1:59*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(7*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(7*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[24*POS_CACHE_WIDTH-1:23*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(7*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(7*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[4*POS_CACHE_WIDTH-1:3*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(7*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(7*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[5*POS_CACHE_WIDTH-1:4*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(8*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(8*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[9*POS_CACHE_WIDTH-1:8*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(8*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(8*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[58*POS_CACHE_WIDTH-1:57*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(8*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(8*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[29*POS_CACHE_WIDTH-1:28*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(8*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(8*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[8*POS_CACHE_WIDTH-1:7*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(8*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(8*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[64*POS_CACHE_WIDTH-1:63*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(8*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(8*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[32*POS_CACHE_WIDTH-1:31*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(8*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(8*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[24*POS_CACHE_WIDTH-1:23*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(8*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(8*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[56*POS_CACHE_WIDTH-1:55*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(8*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(8*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[60*POS_CACHE_WIDTH-1:59*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(8*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(8*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[16*POS_CACHE_WIDTH-1:15*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(8*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(8*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[61*POS_CACHE_WIDTH-1:60*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(8*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(8*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[25*POS_CACHE_WIDTH-1:24*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(8*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(8*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[5*POS_CACHE_WIDTH-1:4*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(8*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(8*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[10*POS_CACHE_WIDTH-1:9*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(9*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(9*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[10*POS_CACHE_WIDTH-1:9*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(9*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(9*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[59*POS_CACHE_WIDTH-1:58*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(9*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(9*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[30*POS_CACHE_WIDTH-1:29*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(9*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(9*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[5*POS_CACHE_WIDTH-1:4*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(9*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(9*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[61*POS_CACHE_WIDTH-1:60*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(9*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(9*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[29*POS_CACHE_WIDTH-1:28*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(9*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(9*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[21*POS_CACHE_WIDTH-1:20*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(9*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(9*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[53*POS_CACHE_WIDTH-1:52*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(9*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(9*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[57*POS_CACHE_WIDTH-1:56*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(9*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(9*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[13*POS_CACHE_WIDTH-1:12*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(9*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(9*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[62*POS_CACHE_WIDTH-1:61*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(9*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(9*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[26*POS_CACHE_WIDTH-1:25*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(9*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(9*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[6*POS_CACHE_WIDTH-1:5*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(9*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(9*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[11*POS_CACHE_WIDTH-1:10*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(10*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(10*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[11*POS_CACHE_WIDTH-1:10*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(10*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(10*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[60*POS_CACHE_WIDTH-1:59*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(10*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(10*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[31*POS_CACHE_WIDTH-1:30*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(10*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(10*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[6*POS_CACHE_WIDTH-1:5*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(10*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(10*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[62*POS_CACHE_WIDTH-1:61*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(10*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(10*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[30*POS_CACHE_WIDTH-1:29*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(10*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(10*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[22*POS_CACHE_WIDTH-1:21*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(10*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(10*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[54*POS_CACHE_WIDTH-1:53*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(10*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(10*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[58*POS_CACHE_WIDTH-1:57*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(10*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(10*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[14*POS_CACHE_WIDTH-1:13*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(10*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(10*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[63*POS_CACHE_WIDTH-1:62*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(10*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(10*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[27*POS_CACHE_WIDTH-1:26*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(10*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(10*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[7*POS_CACHE_WIDTH-1:6*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(10*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(10*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[12*POS_CACHE_WIDTH-1:11*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(11*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(11*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[12*POS_CACHE_WIDTH-1:11*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(11*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(11*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[57*POS_CACHE_WIDTH-1:56*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(11*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(11*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[32*POS_CACHE_WIDTH-1:31*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(11*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(11*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[7*POS_CACHE_WIDTH-1:6*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(11*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(11*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[63*POS_CACHE_WIDTH-1:62*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(11*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(11*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[31*POS_CACHE_WIDTH-1:30*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(11*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(11*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[23*POS_CACHE_WIDTH-1:22*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(11*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(11*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[55*POS_CACHE_WIDTH-1:54*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(11*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(11*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[59*POS_CACHE_WIDTH-1:58*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(11*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(11*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[15*POS_CACHE_WIDTH-1:14*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(11*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(11*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[64*POS_CACHE_WIDTH-1:63*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(11*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(11*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[28*POS_CACHE_WIDTH-1:27*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(11*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(11*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[8*POS_CACHE_WIDTH-1:7*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(11*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(11*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[9*POS_CACHE_WIDTH-1:8*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(12*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(12*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[13*POS_CACHE_WIDTH-1:12*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(12*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(12*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[62*POS_CACHE_WIDTH-1:61*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(12*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(12*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[17*POS_CACHE_WIDTH-1:16*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(12*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(12*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[12*POS_CACHE_WIDTH-1:11*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(12*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(12*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[52*POS_CACHE_WIDTH-1:51*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(12*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(12*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[20*POS_CACHE_WIDTH-1:19*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(12*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(12*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[28*POS_CACHE_WIDTH-1:27*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(12*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(12*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[60*POS_CACHE_WIDTH-1:59*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(12*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(12*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[64*POS_CACHE_WIDTH-1:63*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(12*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(12*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[4*POS_CACHE_WIDTH-1:3*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(12*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(12*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[49*POS_CACHE_WIDTH-1:48*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(12*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(12*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[29*POS_CACHE_WIDTH-1:28*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(12*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(12*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[9*POS_CACHE_WIDTH-1:8*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(12*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(12*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[14*POS_CACHE_WIDTH-1:13*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(13*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(13*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[14*POS_CACHE_WIDTH-1:13*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(13*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(13*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[63*POS_CACHE_WIDTH-1:62*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(13*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(13*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[18*POS_CACHE_WIDTH-1:17*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(13*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(13*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[9*POS_CACHE_WIDTH-1:8*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(13*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(13*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[49*POS_CACHE_WIDTH-1:48*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(13*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(13*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[17*POS_CACHE_WIDTH-1:16*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(13*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(13*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[25*POS_CACHE_WIDTH-1:24*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(13*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(13*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[57*POS_CACHE_WIDTH-1:56*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(13*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(13*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[61*POS_CACHE_WIDTH-1:60*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(13*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(13*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[1*POS_CACHE_WIDTH-1:0*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(13*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(13*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[50*POS_CACHE_WIDTH-1:49*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(13*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(13*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[30*POS_CACHE_WIDTH-1:29*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(13*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(13*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[10*POS_CACHE_WIDTH-1:9*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(13*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(13*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[15*POS_CACHE_WIDTH-1:14*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(14*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(14*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[15*POS_CACHE_WIDTH-1:14*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(14*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(14*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[64*POS_CACHE_WIDTH-1:63*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(14*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(14*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[19*POS_CACHE_WIDTH-1:18*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(14*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(14*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[10*POS_CACHE_WIDTH-1:9*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(14*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(14*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[50*POS_CACHE_WIDTH-1:49*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(14*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(14*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[18*POS_CACHE_WIDTH-1:17*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(14*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(14*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[26*POS_CACHE_WIDTH-1:25*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(14*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(14*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[58*POS_CACHE_WIDTH-1:57*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(14*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(14*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[62*POS_CACHE_WIDTH-1:61*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(14*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(14*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[2*POS_CACHE_WIDTH-1:1*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(14*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(14*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[51*POS_CACHE_WIDTH-1:50*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(14*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(14*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[31*POS_CACHE_WIDTH-1:30*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(14*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(14*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[11*POS_CACHE_WIDTH-1:10*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(14*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(14*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[16*POS_CACHE_WIDTH-1:15*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(15*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(15*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[16*POS_CACHE_WIDTH-1:15*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(15*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(15*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[61*POS_CACHE_WIDTH-1:60*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(15*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(15*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[20*POS_CACHE_WIDTH-1:19*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(15*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(15*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[11*POS_CACHE_WIDTH-1:10*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(15*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(15*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[51*POS_CACHE_WIDTH-1:50*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(15*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(15*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[19*POS_CACHE_WIDTH-1:18*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(15*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(15*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[27*POS_CACHE_WIDTH-1:26*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(15*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(15*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[59*POS_CACHE_WIDTH-1:58*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(15*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(15*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[63*POS_CACHE_WIDTH-1:62*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(15*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(15*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[3*POS_CACHE_WIDTH-1:2*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(15*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(15*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[52*POS_CACHE_WIDTH-1:51*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(15*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(15*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[32*POS_CACHE_WIDTH-1:31*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(15*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(15*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[12*POS_CACHE_WIDTH-1:11*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(15*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(15*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[13*POS_CACHE_WIDTH-1:12*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(16*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(16*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[17*POS_CACHE_WIDTH-1:16*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(16*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(16*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[2*POS_CACHE_WIDTH-1:1*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(16*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(16*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[37*POS_CACHE_WIDTH-1:36*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(16*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(16*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[32*POS_CACHE_WIDTH-1:31*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(16*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(16*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[8*POS_CACHE_WIDTH-1:7*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(16*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(16*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[40*POS_CACHE_WIDTH-1:39*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(16*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(16*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[48*POS_CACHE_WIDTH-1:47*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(16*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(16*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[16*POS_CACHE_WIDTH-1:15*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(16*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(16*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[4*POS_CACHE_WIDTH-1:3*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(16*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(16*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[24*POS_CACHE_WIDTH-1:23*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(16*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(16*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[5*POS_CACHE_WIDTH-1:4*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(16*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(16*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[33*POS_CACHE_WIDTH-1:32*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(16*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(16*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[29*POS_CACHE_WIDTH-1:28*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(16*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(16*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[18*POS_CACHE_WIDTH-1:17*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(17*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(17*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[18*POS_CACHE_WIDTH-1:17*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(17*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(17*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[3*POS_CACHE_WIDTH-1:2*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(17*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(17*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[38*POS_CACHE_WIDTH-1:37*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(17*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(17*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[29*POS_CACHE_WIDTH-1:28*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(17*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(17*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[5*POS_CACHE_WIDTH-1:4*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(17*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(17*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[37*POS_CACHE_WIDTH-1:36*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(17*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(17*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[45*POS_CACHE_WIDTH-1:44*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(17*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(17*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[13*POS_CACHE_WIDTH-1:12*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(17*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(17*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[1*POS_CACHE_WIDTH-1:0*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(17*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(17*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[21*POS_CACHE_WIDTH-1:20*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(17*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(17*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[6*POS_CACHE_WIDTH-1:5*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(17*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(17*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[34*POS_CACHE_WIDTH-1:33*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(17*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(17*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[30*POS_CACHE_WIDTH-1:29*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(17*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(17*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[19*POS_CACHE_WIDTH-1:18*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(18*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(18*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[19*POS_CACHE_WIDTH-1:18*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(18*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(18*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[4*POS_CACHE_WIDTH-1:3*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(18*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(18*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[39*POS_CACHE_WIDTH-1:38*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(18*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(18*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[30*POS_CACHE_WIDTH-1:29*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(18*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(18*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[6*POS_CACHE_WIDTH-1:5*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(18*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(18*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[38*POS_CACHE_WIDTH-1:37*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(18*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(18*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[46*POS_CACHE_WIDTH-1:45*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(18*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(18*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[14*POS_CACHE_WIDTH-1:13*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(18*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(18*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[2*POS_CACHE_WIDTH-1:1*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(18*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(18*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[22*POS_CACHE_WIDTH-1:21*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(18*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(18*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[7*POS_CACHE_WIDTH-1:6*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(18*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(18*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[35*POS_CACHE_WIDTH-1:34*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(18*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(18*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[31*POS_CACHE_WIDTH-1:30*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(18*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(18*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[20*POS_CACHE_WIDTH-1:19*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(19*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(19*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[20*POS_CACHE_WIDTH-1:19*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(19*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(19*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[1*POS_CACHE_WIDTH-1:0*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(19*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(19*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[40*POS_CACHE_WIDTH-1:39*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(19*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(19*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[31*POS_CACHE_WIDTH-1:30*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(19*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(19*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[7*POS_CACHE_WIDTH-1:6*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(19*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(19*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[39*POS_CACHE_WIDTH-1:38*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(19*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(19*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[47*POS_CACHE_WIDTH-1:46*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(19*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(19*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[15*POS_CACHE_WIDTH-1:14*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(19*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(19*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[3*POS_CACHE_WIDTH-1:2*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(19*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(19*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[23*POS_CACHE_WIDTH-1:22*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(19*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(19*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[8*POS_CACHE_WIDTH-1:7*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(19*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(19*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[36*POS_CACHE_WIDTH-1:35*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(19*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(19*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[32*POS_CACHE_WIDTH-1:31*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(19*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(19*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[17*POS_CACHE_WIDTH-1:16*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(20*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(20*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[21*POS_CACHE_WIDTH-1:20*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(20*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(20*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[6*POS_CACHE_WIDTH-1:5*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(20*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(20*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[41*POS_CACHE_WIDTH-1:40*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(20*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(20*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[20*POS_CACHE_WIDTH-1:19*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(20*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(20*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[12*POS_CACHE_WIDTH-1:11*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(20*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(20*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[44*POS_CACHE_WIDTH-1:43*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(20*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(20*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[36*POS_CACHE_WIDTH-1:35*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(20*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(20*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[4*POS_CACHE_WIDTH-1:3*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(20*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(20*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[8*POS_CACHE_WIDTH-1:7*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(20*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(20*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[28*POS_CACHE_WIDTH-1:27*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(20*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(20*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[9*POS_CACHE_WIDTH-1:8*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(20*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(20*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[37*POS_CACHE_WIDTH-1:36*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(20*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(20*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[17*POS_CACHE_WIDTH-1:16*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(20*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(20*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[22*POS_CACHE_WIDTH-1:21*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(21*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(21*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[22*POS_CACHE_WIDTH-1:21*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(21*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(21*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[7*POS_CACHE_WIDTH-1:6*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(21*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(21*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[42*POS_CACHE_WIDTH-1:41*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(21*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(21*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[17*POS_CACHE_WIDTH-1:16*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(21*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(21*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[9*POS_CACHE_WIDTH-1:8*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(21*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(21*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[41*POS_CACHE_WIDTH-1:40*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(21*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(21*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[33*POS_CACHE_WIDTH-1:32*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(21*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(21*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[1*POS_CACHE_WIDTH-1:0*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(21*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(21*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[5*POS_CACHE_WIDTH-1:4*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(21*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(21*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[25*POS_CACHE_WIDTH-1:24*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(21*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(21*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[10*POS_CACHE_WIDTH-1:9*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(21*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(21*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[38*POS_CACHE_WIDTH-1:37*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(21*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(21*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[18*POS_CACHE_WIDTH-1:17*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(21*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(21*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[23*POS_CACHE_WIDTH-1:22*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(22*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(22*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[23*POS_CACHE_WIDTH-1:22*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(22*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(22*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[8*POS_CACHE_WIDTH-1:7*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(22*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(22*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[43*POS_CACHE_WIDTH-1:42*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(22*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(22*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[18*POS_CACHE_WIDTH-1:17*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(22*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(22*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[10*POS_CACHE_WIDTH-1:9*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(22*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(22*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[42*POS_CACHE_WIDTH-1:41*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(22*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(22*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[34*POS_CACHE_WIDTH-1:33*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(22*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(22*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[2*POS_CACHE_WIDTH-1:1*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(22*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(22*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[6*POS_CACHE_WIDTH-1:5*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(22*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(22*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[26*POS_CACHE_WIDTH-1:25*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(22*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(22*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[11*POS_CACHE_WIDTH-1:10*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(22*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(22*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[39*POS_CACHE_WIDTH-1:38*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(22*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(22*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[19*POS_CACHE_WIDTH-1:18*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(22*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(22*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[24*POS_CACHE_WIDTH-1:23*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(23*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(23*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[24*POS_CACHE_WIDTH-1:23*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(23*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(23*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[5*POS_CACHE_WIDTH-1:4*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(23*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(23*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[44*POS_CACHE_WIDTH-1:43*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(23*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(23*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[19*POS_CACHE_WIDTH-1:18*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(23*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(23*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[11*POS_CACHE_WIDTH-1:10*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(23*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(23*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[43*POS_CACHE_WIDTH-1:42*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(23*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(23*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[35*POS_CACHE_WIDTH-1:34*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(23*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(23*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[3*POS_CACHE_WIDTH-1:2*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(23*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(23*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[7*POS_CACHE_WIDTH-1:6*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(23*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(23*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[27*POS_CACHE_WIDTH-1:26*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(23*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(23*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[12*POS_CACHE_WIDTH-1:11*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(23*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(23*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[40*POS_CACHE_WIDTH-1:39*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(23*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(23*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[20*POS_CACHE_WIDTH-1:19*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(23*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(23*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[21*POS_CACHE_WIDTH-1:20*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(24*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(24*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[25*POS_CACHE_WIDTH-1:24*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(24*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(24*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[10*POS_CACHE_WIDTH-1:9*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(24*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(24*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[45*POS_CACHE_WIDTH-1:44*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(24*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(24*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[24*POS_CACHE_WIDTH-1:23*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(24*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(24*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[16*POS_CACHE_WIDTH-1:15*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(24*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(24*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[48*POS_CACHE_WIDTH-1:47*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(24*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(24*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[40*POS_CACHE_WIDTH-1:39*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(24*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(24*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[8*POS_CACHE_WIDTH-1:7*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(24*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(24*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[12*POS_CACHE_WIDTH-1:11*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(24*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(24*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[32*POS_CACHE_WIDTH-1:31*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(24*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(24*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[13*POS_CACHE_WIDTH-1:12*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(24*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(24*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[41*POS_CACHE_WIDTH-1:40*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(24*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(24*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[21*POS_CACHE_WIDTH-1:20*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(24*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(24*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[26*POS_CACHE_WIDTH-1:25*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(25*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(25*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[26*POS_CACHE_WIDTH-1:25*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(25*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(25*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[11*POS_CACHE_WIDTH-1:10*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(25*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(25*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[46*POS_CACHE_WIDTH-1:45*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(25*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(25*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[21*POS_CACHE_WIDTH-1:20*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(25*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(25*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[13*POS_CACHE_WIDTH-1:12*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(25*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(25*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[45*POS_CACHE_WIDTH-1:44*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(25*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(25*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[37*POS_CACHE_WIDTH-1:36*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(25*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(25*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[5*POS_CACHE_WIDTH-1:4*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(25*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(25*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[9*POS_CACHE_WIDTH-1:8*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(25*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(25*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[29*POS_CACHE_WIDTH-1:28*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(25*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(25*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[14*POS_CACHE_WIDTH-1:13*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(25*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(25*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[42*POS_CACHE_WIDTH-1:41*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(25*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(25*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[22*POS_CACHE_WIDTH-1:21*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(25*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(25*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[27*POS_CACHE_WIDTH-1:26*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(26*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(26*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[27*POS_CACHE_WIDTH-1:26*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(26*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(26*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[12*POS_CACHE_WIDTH-1:11*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(26*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(26*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[47*POS_CACHE_WIDTH-1:46*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(26*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(26*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[22*POS_CACHE_WIDTH-1:21*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(26*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(26*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[14*POS_CACHE_WIDTH-1:13*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(26*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(26*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[46*POS_CACHE_WIDTH-1:45*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(26*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(26*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[38*POS_CACHE_WIDTH-1:37*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(26*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(26*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[6*POS_CACHE_WIDTH-1:5*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(26*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(26*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[10*POS_CACHE_WIDTH-1:9*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(26*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(26*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[30*POS_CACHE_WIDTH-1:29*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(26*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(26*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[15*POS_CACHE_WIDTH-1:14*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(26*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(26*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[43*POS_CACHE_WIDTH-1:42*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(26*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(26*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[23*POS_CACHE_WIDTH-1:22*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(26*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(26*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[28*POS_CACHE_WIDTH-1:27*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(27*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(27*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[28*POS_CACHE_WIDTH-1:27*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(27*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(27*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[9*POS_CACHE_WIDTH-1:8*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(27*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(27*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[48*POS_CACHE_WIDTH-1:47*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(27*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(27*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[23*POS_CACHE_WIDTH-1:22*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(27*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(27*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[15*POS_CACHE_WIDTH-1:14*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(27*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(27*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[47*POS_CACHE_WIDTH-1:46*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(27*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(27*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[39*POS_CACHE_WIDTH-1:38*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(27*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(27*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[7*POS_CACHE_WIDTH-1:6*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(27*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(27*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[11*POS_CACHE_WIDTH-1:10*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(27*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(27*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[31*POS_CACHE_WIDTH-1:30*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(27*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(27*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[16*POS_CACHE_WIDTH-1:15*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(27*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(27*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[44*POS_CACHE_WIDTH-1:43*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(27*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(27*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[24*POS_CACHE_WIDTH-1:23*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(27*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(27*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[25*POS_CACHE_WIDTH-1:24*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(28*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(28*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[29*POS_CACHE_WIDTH-1:28*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(28*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(28*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[14*POS_CACHE_WIDTH-1:13*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(28*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(28*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[33*POS_CACHE_WIDTH-1:32*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(28*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(28*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[28*POS_CACHE_WIDTH-1:27*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(28*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(28*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[4*POS_CACHE_WIDTH-1:3*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(28*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(28*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[36*POS_CACHE_WIDTH-1:35*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(28*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(28*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[44*POS_CACHE_WIDTH-1:43*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(28*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(28*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[12*POS_CACHE_WIDTH-1:11*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(28*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(28*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[16*POS_CACHE_WIDTH-1:15*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(28*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(28*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[20*POS_CACHE_WIDTH-1:19*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(28*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(28*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[1*POS_CACHE_WIDTH-1:0*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(28*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(28*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[45*POS_CACHE_WIDTH-1:44*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(28*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(28*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[25*POS_CACHE_WIDTH-1:24*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(28*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(28*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[30*POS_CACHE_WIDTH-1:29*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(29*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(29*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[30*POS_CACHE_WIDTH-1:29*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(29*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(29*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[15*POS_CACHE_WIDTH-1:14*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(29*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(29*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[34*POS_CACHE_WIDTH-1:33*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(29*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(29*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[25*POS_CACHE_WIDTH-1:24*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(29*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(29*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[1*POS_CACHE_WIDTH-1:0*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(29*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(29*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[33*POS_CACHE_WIDTH-1:32*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(29*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(29*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[41*POS_CACHE_WIDTH-1:40*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(29*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(29*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[9*POS_CACHE_WIDTH-1:8*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(29*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(29*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[13*POS_CACHE_WIDTH-1:12*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(29*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(29*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[17*POS_CACHE_WIDTH-1:16*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(29*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(29*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[2*POS_CACHE_WIDTH-1:1*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(29*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(29*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[46*POS_CACHE_WIDTH-1:45*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(29*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(29*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[26*POS_CACHE_WIDTH-1:25*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(29*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(29*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[31*POS_CACHE_WIDTH-1:30*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(30*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(30*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[31*POS_CACHE_WIDTH-1:30*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(30*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(30*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[16*POS_CACHE_WIDTH-1:15*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(30*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(30*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[35*POS_CACHE_WIDTH-1:34*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(30*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(30*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[26*POS_CACHE_WIDTH-1:25*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(30*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(30*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[2*POS_CACHE_WIDTH-1:1*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(30*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(30*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[34*POS_CACHE_WIDTH-1:33*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(30*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(30*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[42*POS_CACHE_WIDTH-1:41*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(30*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(30*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[10*POS_CACHE_WIDTH-1:9*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(30*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(30*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[14*POS_CACHE_WIDTH-1:13*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(30*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(30*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[18*POS_CACHE_WIDTH-1:17*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(30*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(30*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[3*POS_CACHE_WIDTH-1:2*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(30*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(30*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[47*POS_CACHE_WIDTH-1:46*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(30*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(30*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[27*POS_CACHE_WIDTH-1:26*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(30*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(30*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[32*POS_CACHE_WIDTH-1:31*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(31*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(31*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[32*POS_CACHE_WIDTH-1:31*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(31*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(31*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[13*POS_CACHE_WIDTH-1:12*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(31*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(31*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[36*POS_CACHE_WIDTH-1:35*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(31*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(31*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[27*POS_CACHE_WIDTH-1:26*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(31*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(31*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[3*POS_CACHE_WIDTH-1:2*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(31*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(31*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[35*POS_CACHE_WIDTH-1:34*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(31*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(31*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[43*POS_CACHE_WIDTH-1:42*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(31*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(31*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[11*POS_CACHE_WIDTH-1:10*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(31*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(31*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[15*POS_CACHE_WIDTH-1:14*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(31*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(31*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[19*POS_CACHE_WIDTH-1:18*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(31*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(31*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[4*POS_CACHE_WIDTH-1:3*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(31*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(31*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[48*POS_CACHE_WIDTH-1:47*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(31*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(31*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[28*POS_CACHE_WIDTH-1:27*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(31*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(31*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[29*POS_CACHE_WIDTH-1:28*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(32*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(32*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[33*POS_CACHE_WIDTH-1:32*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(32*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(32*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[18*POS_CACHE_WIDTH-1:17*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(32*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(32*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[53*POS_CACHE_WIDTH-1:52*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(32*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(32*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[48*POS_CACHE_WIDTH-1:47*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(32*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(32*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[24*POS_CACHE_WIDTH-1:23*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(32*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(32*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[56*POS_CACHE_WIDTH-1:55*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(32*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(32*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[64*POS_CACHE_WIDTH-1:63*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(32*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(32*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[32*POS_CACHE_WIDTH-1:31*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(32*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(32*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[20*POS_CACHE_WIDTH-1:19*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(32*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(32*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[40*POS_CACHE_WIDTH-1:39*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(32*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(32*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[21*POS_CACHE_WIDTH-1:20*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(32*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(32*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[49*POS_CACHE_WIDTH-1:48*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(32*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(32*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[45*POS_CACHE_WIDTH-1:44*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(32*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(32*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[34*POS_CACHE_WIDTH-1:33*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(33*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(33*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[34*POS_CACHE_WIDTH-1:33*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(33*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(33*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[19*POS_CACHE_WIDTH-1:18*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(33*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(33*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[54*POS_CACHE_WIDTH-1:53*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(33*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(33*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[45*POS_CACHE_WIDTH-1:44*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(33*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(33*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[21*POS_CACHE_WIDTH-1:20*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(33*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(33*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[53*POS_CACHE_WIDTH-1:52*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(33*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(33*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[61*POS_CACHE_WIDTH-1:60*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(33*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(33*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[29*POS_CACHE_WIDTH-1:28*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(33*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(33*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[17*POS_CACHE_WIDTH-1:16*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(33*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(33*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[37*POS_CACHE_WIDTH-1:36*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(33*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(33*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[22*POS_CACHE_WIDTH-1:21*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(33*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(33*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[50*POS_CACHE_WIDTH-1:49*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(33*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(33*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[46*POS_CACHE_WIDTH-1:45*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(33*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(33*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[35*POS_CACHE_WIDTH-1:34*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(34*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(34*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[35*POS_CACHE_WIDTH-1:34*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(34*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(34*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[20*POS_CACHE_WIDTH-1:19*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(34*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(34*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[55*POS_CACHE_WIDTH-1:54*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(34*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(34*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[46*POS_CACHE_WIDTH-1:45*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(34*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(34*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[22*POS_CACHE_WIDTH-1:21*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(34*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(34*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[54*POS_CACHE_WIDTH-1:53*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(34*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(34*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[62*POS_CACHE_WIDTH-1:61*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(34*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(34*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[30*POS_CACHE_WIDTH-1:29*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(34*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(34*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[18*POS_CACHE_WIDTH-1:17*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(34*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(34*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[38*POS_CACHE_WIDTH-1:37*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(34*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(34*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[23*POS_CACHE_WIDTH-1:22*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(34*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(34*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[51*POS_CACHE_WIDTH-1:50*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(34*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(34*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[47*POS_CACHE_WIDTH-1:46*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(34*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(34*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[36*POS_CACHE_WIDTH-1:35*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(35*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(35*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[36*POS_CACHE_WIDTH-1:35*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(35*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(35*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[17*POS_CACHE_WIDTH-1:16*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(35*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(35*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[56*POS_CACHE_WIDTH-1:55*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(35*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(35*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[47*POS_CACHE_WIDTH-1:46*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(35*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(35*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[23*POS_CACHE_WIDTH-1:22*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(35*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(35*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[55*POS_CACHE_WIDTH-1:54*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(35*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(35*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[63*POS_CACHE_WIDTH-1:62*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(35*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(35*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[31*POS_CACHE_WIDTH-1:30*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(35*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(35*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[19*POS_CACHE_WIDTH-1:18*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(35*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(35*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[39*POS_CACHE_WIDTH-1:38*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(35*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(35*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[24*POS_CACHE_WIDTH-1:23*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(35*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(35*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[52*POS_CACHE_WIDTH-1:51*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(35*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(35*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[48*POS_CACHE_WIDTH-1:47*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(35*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(35*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[33*POS_CACHE_WIDTH-1:32*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(36*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(36*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[37*POS_CACHE_WIDTH-1:36*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(36*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(36*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[22*POS_CACHE_WIDTH-1:21*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(36*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(36*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[57*POS_CACHE_WIDTH-1:56*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(36*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(36*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[36*POS_CACHE_WIDTH-1:35*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(36*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(36*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[28*POS_CACHE_WIDTH-1:27*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(36*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(36*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[60*POS_CACHE_WIDTH-1:59*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(36*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(36*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[52*POS_CACHE_WIDTH-1:51*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(36*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(36*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[20*POS_CACHE_WIDTH-1:19*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(36*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(36*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[24*POS_CACHE_WIDTH-1:23*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(36*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(36*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[44*POS_CACHE_WIDTH-1:43*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(36*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(36*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[25*POS_CACHE_WIDTH-1:24*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(36*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(36*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[53*POS_CACHE_WIDTH-1:52*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(36*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(36*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[33*POS_CACHE_WIDTH-1:32*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(36*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(36*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[38*POS_CACHE_WIDTH-1:37*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(37*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(37*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[38*POS_CACHE_WIDTH-1:37*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(37*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(37*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[23*POS_CACHE_WIDTH-1:22*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(37*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(37*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[58*POS_CACHE_WIDTH-1:57*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(37*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(37*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[33*POS_CACHE_WIDTH-1:32*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(37*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(37*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[25*POS_CACHE_WIDTH-1:24*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(37*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(37*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[57*POS_CACHE_WIDTH-1:56*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(37*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(37*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[49*POS_CACHE_WIDTH-1:48*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(37*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(37*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[17*POS_CACHE_WIDTH-1:16*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(37*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(37*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[21*POS_CACHE_WIDTH-1:20*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(37*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(37*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[41*POS_CACHE_WIDTH-1:40*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(37*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(37*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[26*POS_CACHE_WIDTH-1:25*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(37*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(37*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[54*POS_CACHE_WIDTH-1:53*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(37*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(37*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[34*POS_CACHE_WIDTH-1:33*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(37*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(37*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[39*POS_CACHE_WIDTH-1:38*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(38*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(38*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[39*POS_CACHE_WIDTH-1:38*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(38*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(38*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[24*POS_CACHE_WIDTH-1:23*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(38*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(38*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[59*POS_CACHE_WIDTH-1:58*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(38*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(38*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[34*POS_CACHE_WIDTH-1:33*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(38*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(38*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[26*POS_CACHE_WIDTH-1:25*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(38*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(38*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[58*POS_CACHE_WIDTH-1:57*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(38*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(38*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[50*POS_CACHE_WIDTH-1:49*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(38*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(38*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[18*POS_CACHE_WIDTH-1:17*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(38*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(38*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[22*POS_CACHE_WIDTH-1:21*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(38*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(38*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[42*POS_CACHE_WIDTH-1:41*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(38*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(38*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[27*POS_CACHE_WIDTH-1:26*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(38*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(38*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[55*POS_CACHE_WIDTH-1:54*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(38*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(38*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[35*POS_CACHE_WIDTH-1:34*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(38*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(38*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[40*POS_CACHE_WIDTH-1:39*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(39*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(39*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[40*POS_CACHE_WIDTH-1:39*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(39*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(39*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[21*POS_CACHE_WIDTH-1:20*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(39*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(39*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[60*POS_CACHE_WIDTH-1:59*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(39*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(39*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[35*POS_CACHE_WIDTH-1:34*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(39*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(39*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[27*POS_CACHE_WIDTH-1:26*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(39*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(39*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[59*POS_CACHE_WIDTH-1:58*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(39*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(39*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[51*POS_CACHE_WIDTH-1:50*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(39*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(39*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[19*POS_CACHE_WIDTH-1:18*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(39*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(39*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[23*POS_CACHE_WIDTH-1:22*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(39*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(39*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[43*POS_CACHE_WIDTH-1:42*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(39*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(39*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[28*POS_CACHE_WIDTH-1:27*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(39*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(39*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[56*POS_CACHE_WIDTH-1:55*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(39*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(39*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[36*POS_CACHE_WIDTH-1:35*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(39*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(39*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[37*POS_CACHE_WIDTH-1:36*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(40*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(40*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[41*POS_CACHE_WIDTH-1:40*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(40*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(40*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[26*POS_CACHE_WIDTH-1:25*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(40*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(40*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[61*POS_CACHE_WIDTH-1:60*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(40*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(40*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[40*POS_CACHE_WIDTH-1:39*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(40*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(40*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[32*POS_CACHE_WIDTH-1:31*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(40*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(40*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[64*POS_CACHE_WIDTH-1:63*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(40*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(40*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[56*POS_CACHE_WIDTH-1:55*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(40*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(40*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[24*POS_CACHE_WIDTH-1:23*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(40*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(40*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[28*POS_CACHE_WIDTH-1:27*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(40*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(40*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[48*POS_CACHE_WIDTH-1:47*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(40*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(40*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[29*POS_CACHE_WIDTH-1:28*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(40*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(40*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[57*POS_CACHE_WIDTH-1:56*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(40*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(40*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[37*POS_CACHE_WIDTH-1:36*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(40*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(40*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[42*POS_CACHE_WIDTH-1:41*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(41*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(41*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[42*POS_CACHE_WIDTH-1:41*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(41*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(41*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[27*POS_CACHE_WIDTH-1:26*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(41*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(41*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[62*POS_CACHE_WIDTH-1:61*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(41*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(41*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[37*POS_CACHE_WIDTH-1:36*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(41*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(41*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[29*POS_CACHE_WIDTH-1:28*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(41*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(41*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[61*POS_CACHE_WIDTH-1:60*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(41*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(41*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[53*POS_CACHE_WIDTH-1:52*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(41*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(41*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[21*POS_CACHE_WIDTH-1:20*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(41*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(41*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[25*POS_CACHE_WIDTH-1:24*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(41*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(41*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[45*POS_CACHE_WIDTH-1:44*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(41*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(41*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[30*POS_CACHE_WIDTH-1:29*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(41*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(41*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[58*POS_CACHE_WIDTH-1:57*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(41*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(41*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[38*POS_CACHE_WIDTH-1:37*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(41*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(41*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[43*POS_CACHE_WIDTH-1:42*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(42*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(42*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[43*POS_CACHE_WIDTH-1:42*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(42*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(42*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[28*POS_CACHE_WIDTH-1:27*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(42*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(42*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[63*POS_CACHE_WIDTH-1:62*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(42*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(42*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[38*POS_CACHE_WIDTH-1:37*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(42*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(42*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[30*POS_CACHE_WIDTH-1:29*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(42*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(42*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[62*POS_CACHE_WIDTH-1:61*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(42*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(42*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[54*POS_CACHE_WIDTH-1:53*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(42*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(42*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[22*POS_CACHE_WIDTH-1:21*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(42*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(42*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[26*POS_CACHE_WIDTH-1:25*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(42*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(42*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[46*POS_CACHE_WIDTH-1:45*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(42*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(42*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[31*POS_CACHE_WIDTH-1:30*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(42*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(42*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[59*POS_CACHE_WIDTH-1:58*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(42*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(42*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[39*POS_CACHE_WIDTH-1:38*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(42*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(42*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[44*POS_CACHE_WIDTH-1:43*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(43*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(43*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[44*POS_CACHE_WIDTH-1:43*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(43*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(43*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[25*POS_CACHE_WIDTH-1:24*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(43*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(43*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[64*POS_CACHE_WIDTH-1:63*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(43*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(43*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[39*POS_CACHE_WIDTH-1:38*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(43*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(43*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[31*POS_CACHE_WIDTH-1:30*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(43*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(43*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[63*POS_CACHE_WIDTH-1:62*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(43*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(43*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[55*POS_CACHE_WIDTH-1:54*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(43*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(43*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[23*POS_CACHE_WIDTH-1:22*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(43*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(43*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[27*POS_CACHE_WIDTH-1:26*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(43*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(43*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[47*POS_CACHE_WIDTH-1:46*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(43*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(43*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[32*POS_CACHE_WIDTH-1:31*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(43*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(43*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[60*POS_CACHE_WIDTH-1:59*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(43*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(43*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[40*POS_CACHE_WIDTH-1:39*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(43*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(43*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[41*POS_CACHE_WIDTH-1:40*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(44*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(44*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[45*POS_CACHE_WIDTH-1:44*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(44*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(44*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[30*POS_CACHE_WIDTH-1:29*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(44*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(44*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[49*POS_CACHE_WIDTH-1:48*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(44*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(44*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[44*POS_CACHE_WIDTH-1:43*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(44*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(44*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[20*POS_CACHE_WIDTH-1:19*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(44*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(44*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[52*POS_CACHE_WIDTH-1:51*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(44*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(44*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[60*POS_CACHE_WIDTH-1:59*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(44*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(44*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[28*POS_CACHE_WIDTH-1:27*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(44*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(44*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[32*POS_CACHE_WIDTH-1:31*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(44*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(44*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[36*POS_CACHE_WIDTH-1:35*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(44*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(44*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[17*POS_CACHE_WIDTH-1:16*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(44*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(44*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[61*POS_CACHE_WIDTH-1:60*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(44*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(44*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[41*POS_CACHE_WIDTH-1:40*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(44*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(44*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[46*POS_CACHE_WIDTH-1:45*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(45*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(45*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[46*POS_CACHE_WIDTH-1:45*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(45*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(45*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[31*POS_CACHE_WIDTH-1:30*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(45*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(45*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[50*POS_CACHE_WIDTH-1:49*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(45*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(45*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[41*POS_CACHE_WIDTH-1:40*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(45*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(45*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[17*POS_CACHE_WIDTH-1:16*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(45*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(45*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[49*POS_CACHE_WIDTH-1:48*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(45*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(45*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[57*POS_CACHE_WIDTH-1:56*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(45*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(45*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[25*POS_CACHE_WIDTH-1:24*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(45*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(45*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[29*POS_CACHE_WIDTH-1:28*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(45*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(45*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[33*POS_CACHE_WIDTH-1:32*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(45*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(45*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[18*POS_CACHE_WIDTH-1:17*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(45*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(45*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[62*POS_CACHE_WIDTH-1:61*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(45*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(45*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[42*POS_CACHE_WIDTH-1:41*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(45*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(45*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[47*POS_CACHE_WIDTH-1:46*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(46*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(46*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[47*POS_CACHE_WIDTH-1:46*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(46*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(46*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[32*POS_CACHE_WIDTH-1:31*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(46*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(46*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[51*POS_CACHE_WIDTH-1:50*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(46*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(46*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[42*POS_CACHE_WIDTH-1:41*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(46*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(46*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[18*POS_CACHE_WIDTH-1:17*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(46*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(46*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[50*POS_CACHE_WIDTH-1:49*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(46*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(46*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[58*POS_CACHE_WIDTH-1:57*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(46*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(46*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[26*POS_CACHE_WIDTH-1:25*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(46*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(46*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[30*POS_CACHE_WIDTH-1:29*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(46*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(46*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[34*POS_CACHE_WIDTH-1:33*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(46*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(46*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[19*POS_CACHE_WIDTH-1:18*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(46*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(46*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[63*POS_CACHE_WIDTH-1:62*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(46*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(46*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[43*POS_CACHE_WIDTH-1:42*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(46*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(46*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[48*POS_CACHE_WIDTH-1:47*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(47*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(47*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[48*POS_CACHE_WIDTH-1:47*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(47*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(47*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[29*POS_CACHE_WIDTH-1:28*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(47*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(47*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[52*POS_CACHE_WIDTH-1:51*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(47*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(47*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[43*POS_CACHE_WIDTH-1:42*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(47*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(47*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[19*POS_CACHE_WIDTH-1:18*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(47*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(47*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[51*POS_CACHE_WIDTH-1:50*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(47*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(47*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[59*POS_CACHE_WIDTH-1:58*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(47*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(47*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[27*POS_CACHE_WIDTH-1:26*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(47*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(47*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[31*POS_CACHE_WIDTH-1:30*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(47*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(47*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[35*POS_CACHE_WIDTH-1:34*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(47*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(47*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[20*POS_CACHE_WIDTH-1:19*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(47*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(47*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[64*POS_CACHE_WIDTH-1:63*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(47*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(47*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[44*POS_CACHE_WIDTH-1:43*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(47*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(47*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[45*POS_CACHE_WIDTH-1:44*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(48*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(48*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[49*POS_CACHE_WIDTH-1:48*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(48*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(48*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[34*POS_CACHE_WIDTH-1:33*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(48*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(48*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[5*POS_CACHE_WIDTH-1:4*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(48*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(48*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[64*POS_CACHE_WIDTH-1:63*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(48*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(48*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[40*POS_CACHE_WIDTH-1:39*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(48*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(48*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[8*POS_CACHE_WIDTH-1:7*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(48*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(48*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[16*POS_CACHE_WIDTH-1:15*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(48*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(48*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[48*POS_CACHE_WIDTH-1:47*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(48*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(48*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[36*POS_CACHE_WIDTH-1:35*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(48*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(48*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[56*POS_CACHE_WIDTH-1:55*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(48*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(48*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[37*POS_CACHE_WIDTH-1:36*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(48*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(48*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[1*POS_CACHE_WIDTH-1:0*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(48*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(48*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[61*POS_CACHE_WIDTH-1:60*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(48*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(48*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[50*POS_CACHE_WIDTH-1:49*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(49*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(49*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[50*POS_CACHE_WIDTH-1:49*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(49*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(49*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[35*POS_CACHE_WIDTH-1:34*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(49*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(49*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[6*POS_CACHE_WIDTH-1:5*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(49*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(49*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[61*POS_CACHE_WIDTH-1:60*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(49*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(49*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[37*POS_CACHE_WIDTH-1:36*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(49*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(49*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[5*POS_CACHE_WIDTH-1:4*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(49*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(49*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[13*POS_CACHE_WIDTH-1:12*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(49*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(49*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[45*POS_CACHE_WIDTH-1:44*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(49*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(49*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[33*POS_CACHE_WIDTH-1:32*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(49*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(49*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[53*POS_CACHE_WIDTH-1:52*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(49*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(49*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[38*POS_CACHE_WIDTH-1:37*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(49*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(49*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[2*POS_CACHE_WIDTH-1:1*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(49*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(49*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[62*POS_CACHE_WIDTH-1:61*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(49*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(49*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[51*POS_CACHE_WIDTH-1:50*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(50*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(50*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[51*POS_CACHE_WIDTH-1:50*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(50*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(50*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[36*POS_CACHE_WIDTH-1:35*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(50*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(50*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[7*POS_CACHE_WIDTH-1:6*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(50*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(50*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[62*POS_CACHE_WIDTH-1:61*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(50*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(50*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[38*POS_CACHE_WIDTH-1:37*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(50*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(50*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[6*POS_CACHE_WIDTH-1:5*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(50*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(50*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[14*POS_CACHE_WIDTH-1:13*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(50*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(50*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[46*POS_CACHE_WIDTH-1:45*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(50*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(50*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[34*POS_CACHE_WIDTH-1:33*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(50*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(50*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[54*POS_CACHE_WIDTH-1:53*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(50*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(50*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[39*POS_CACHE_WIDTH-1:38*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(50*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(50*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[3*POS_CACHE_WIDTH-1:2*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(50*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(50*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[63*POS_CACHE_WIDTH-1:62*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(50*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(50*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[52*POS_CACHE_WIDTH-1:51*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(51*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(51*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[52*POS_CACHE_WIDTH-1:51*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(51*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(51*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[33*POS_CACHE_WIDTH-1:32*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(51*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(51*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[8*POS_CACHE_WIDTH-1:7*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(51*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(51*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[63*POS_CACHE_WIDTH-1:62*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(51*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(51*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[39*POS_CACHE_WIDTH-1:38*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(51*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(51*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[7*POS_CACHE_WIDTH-1:6*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(51*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(51*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[15*POS_CACHE_WIDTH-1:14*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(51*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(51*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[47*POS_CACHE_WIDTH-1:46*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(51*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(51*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[35*POS_CACHE_WIDTH-1:34*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(51*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(51*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[55*POS_CACHE_WIDTH-1:54*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(51*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(51*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[40*POS_CACHE_WIDTH-1:39*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(51*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(51*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[4*POS_CACHE_WIDTH-1:3*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(51*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(51*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[64*POS_CACHE_WIDTH-1:63*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(51*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(51*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[49*POS_CACHE_WIDTH-1:48*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(52*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(52*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[53*POS_CACHE_WIDTH-1:52*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(52*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(52*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[38*POS_CACHE_WIDTH-1:37*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(52*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(52*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[9*POS_CACHE_WIDTH-1:8*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(52*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(52*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[52*POS_CACHE_WIDTH-1:51*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(52*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(52*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[44*POS_CACHE_WIDTH-1:43*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(52*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(52*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[12*POS_CACHE_WIDTH-1:11*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(52*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(52*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[4*POS_CACHE_WIDTH-1:3*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(52*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(52*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[36*POS_CACHE_WIDTH-1:35*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(52*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(52*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[40*POS_CACHE_WIDTH-1:39*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(52*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(52*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[60*POS_CACHE_WIDTH-1:59*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(52*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(52*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[41*POS_CACHE_WIDTH-1:40*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(52*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(52*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[5*POS_CACHE_WIDTH-1:4*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(52*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(52*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[49*POS_CACHE_WIDTH-1:48*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(52*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(52*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[54*POS_CACHE_WIDTH-1:53*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(53*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(53*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[54*POS_CACHE_WIDTH-1:53*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(53*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(53*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[39*POS_CACHE_WIDTH-1:38*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(53*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(53*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[10*POS_CACHE_WIDTH-1:9*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(53*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(53*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[49*POS_CACHE_WIDTH-1:48*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(53*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(53*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[41*POS_CACHE_WIDTH-1:40*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(53*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(53*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[9*POS_CACHE_WIDTH-1:8*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(53*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(53*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[1*POS_CACHE_WIDTH-1:0*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(53*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(53*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[33*POS_CACHE_WIDTH-1:32*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(53*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(53*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[37*POS_CACHE_WIDTH-1:36*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(53*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(53*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[57*POS_CACHE_WIDTH-1:56*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(53*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(53*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[42*POS_CACHE_WIDTH-1:41*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(53*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(53*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[6*POS_CACHE_WIDTH-1:5*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(53*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(53*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[50*POS_CACHE_WIDTH-1:49*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(53*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(53*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[55*POS_CACHE_WIDTH-1:54*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(54*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(54*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[55*POS_CACHE_WIDTH-1:54*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(54*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(54*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[40*POS_CACHE_WIDTH-1:39*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(54*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(54*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[11*POS_CACHE_WIDTH-1:10*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(54*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(54*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[50*POS_CACHE_WIDTH-1:49*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(54*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(54*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[42*POS_CACHE_WIDTH-1:41*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(54*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(54*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[10*POS_CACHE_WIDTH-1:9*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(54*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(54*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[2*POS_CACHE_WIDTH-1:1*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(54*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(54*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[34*POS_CACHE_WIDTH-1:33*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(54*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(54*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[38*POS_CACHE_WIDTH-1:37*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(54*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(54*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[58*POS_CACHE_WIDTH-1:57*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(54*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(54*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[43*POS_CACHE_WIDTH-1:42*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(54*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(54*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[7*POS_CACHE_WIDTH-1:6*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(54*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(54*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[51*POS_CACHE_WIDTH-1:50*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(54*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(54*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[56*POS_CACHE_WIDTH-1:55*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(55*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(55*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[56*POS_CACHE_WIDTH-1:55*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(55*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(55*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[37*POS_CACHE_WIDTH-1:36*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(55*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(55*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[12*POS_CACHE_WIDTH-1:11*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(55*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(55*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[51*POS_CACHE_WIDTH-1:50*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(55*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(55*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[43*POS_CACHE_WIDTH-1:42*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(55*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(55*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[11*POS_CACHE_WIDTH-1:10*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(55*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(55*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[3*POS_CACHE_WIDTH-1:2*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(55*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(55*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[35*POS_CACHE_WIDTH-1:34*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(55*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(55*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[39*POS_CACHE_WIDTH-1:38*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(55*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(55*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[59*POS_CACHE_WIDTH-1:58*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(55*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(55*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[44*POS_CACHE_WIDTH-1:43*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(55*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(55*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[8*POS_CACHE_WIDTH-1:7*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(55*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(55*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[52*POS_CACHE_WIDTH-1:51*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(55*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(55*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[53*POS_CACHE_WIDTH-1:52*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(56*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(56*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[57*POS_CACHE_WIDTH-1:56*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(56*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(56*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[42*POS_CACHE_WIDTH-1:41*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(56*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(56*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[13*POS_CACHE_WIDTH-1:12*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(56*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(56*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[56*POS_CACHE_WIDTH-1:55*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(56*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(56*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[48*POS_CACHE_WIDTH-1:47*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(56*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(56*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[16*POS_CACHE_WIDTH-1:15*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(56*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(56*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[8*POS_CACHE_WIDTH-1:7*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(56*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(56*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[40*POS_CACHE_WIDTH-1:39*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(56*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(56*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[44*POS_CACHE_WIDTH-1:43*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(56*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(56*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[64*POS_CACHE_WIDTH-1:63*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(56*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(56*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[45*POS_CACHE_WIDTH-1:44*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(56*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(56*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[9*POS_CACHE_WIDTH-1:8*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(56*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(56*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[53*POS_CACHE_WIDTH-1:52*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(56*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(56*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[58*POS_CACHE_WIDTH-1:57*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(57*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(57*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[58*POS_CACHE_WIDTH-1:57*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(57*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(57*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[43*POS_CACHE_WIDTH-1:42*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(57*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(57*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[14*POS_CACHE_WIDTH-1:13*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(57*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(57*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[53*POS_CACHE_WIDTH-1:52*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(57*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(57*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[45*POS_CACHE_WIDTH-1:44*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(57*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(57*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[13*POS_CACHE_WIDTH-1:12*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(57*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(57*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[5*POS_CACHE_WIDTH-1:4*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(57*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(57*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[37*POS_CACHE_WIDTH-1:36*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(57*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(57*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[41*POS_CACHE_WIDTH-1:40*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(57*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(57*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[61*POS_CACHE_WIDTH-1:60*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(57*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(57*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[46*POS_CACHE_WIDTH-1:45*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(57*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(57*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[10*POS_CACHE_WIDTH-1:9*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(57*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(57*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[54*POS_CACHE_WIDTH-1:53*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(57*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(57*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[59*POS_CACHE_WIDTH-1:58*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(58*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(58*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[59*POS_CACHE_WIDTH-1:58*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(58*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(58*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[44*POS_CACHE_WIDTH-1:43*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(58*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(58*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[15*POS_CACHE_WIDTH-1:14*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(58*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(58*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[54*POS_CACHE_WIDTH-1:53*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(58*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(58*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[46*POS_CACHE_WIDTH-1:45*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(58*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(58*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[14*POS_CACHE_WIDTH-1:13*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(58*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(58*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[6*POS_CACHE_WIDTH-1:5*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(58*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(58*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[38*POS_CACHE_WIDTH-1:37*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(58*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(58*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[42*POS_CACHE_WIDTH-1:41*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(58*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(58*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[62*POS_CACHE_WIDTH-1:61*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(58*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(58*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[47*POS_CACHE_WIDTH-1:46*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(58*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(58*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[11*POS_CACHE_WIDTH-1:10*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(58*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(58*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[55*POS_CACHE_WIDTH-1:54*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(58*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(58*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[60*POS_CACHE_WIDTH-1:59*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(59*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(59*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[60*POS_CACHE_WIDTH-1:59*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(59*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(59*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[41*POS_CACHE_WIDTH-1:40*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(59*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(59*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[16*POS_CACHE_WIDTH-1:15*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(59*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(59*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[55*POS_CACHE_WIDTH-1:54*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(59*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(59*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[47*POS_CACHE_WIDTH-1:46*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(59*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(59*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[15*POS_CACHE_WIDTH-1:14*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(59*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(59*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[7*POS_CACHE_WIDTH-1:6*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(59*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(59*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[39*POS_CACHE_WIDTH-1:38*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(59*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(59*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[43*POS_CACHE_WIDTH-1:42*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(59*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(59*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[63*POS_CACHE_WIDTH-1:62*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(59*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(59*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[48*POS_CACHE_WIDTH-1:47*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(59*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(59*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[12*POS_CACHE_WIDTH-1:11*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(59*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(59*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[56*POS_CACHE_WIDTH-1:55*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(59*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(59*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[57*POS_CACHE_WIDTH-1:56*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(60*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(60*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[61*POS_CACHE_WIDTH-1:60*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(60*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(60*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[46*POS_CACHE_WIDTH-1:45*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(60*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(60*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[1*POS_CACHE_WIDTH-1:0*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(60*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(60*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[60*POS_CACHE_WIDTH-1:59*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(60*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(60*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[36*POS_CACHE_WIDTH-1:35*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(60*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(60*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[4*POS_CACHE_WIDTH-1:3*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(60*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(60*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[12*POS_CACHE_WIDTH-1:11*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(60*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(60*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[44*POS_CACHE_WIDTH-1:43*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(60*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(60*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[48*POS_CACHE_WIDTH-1:47*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(60*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(60*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[52*POS_CACHE_WIDTH-1:51*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(60*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(60*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[33*POS_CACHE_WIDTH-1:32*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(60*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(60*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[13*POS_CACHE_WIDTH-1:12*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(60*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(60*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[57*POS_CACHE_WIDTH-1:56*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(60*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(60*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[62*POS_CACHE_WIDTH-1:61*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(61*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(61*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[62*POS_CACHE_WIDTH-1:61*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(61*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(61*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[47*POS_CACHE_WIDTH-1:46*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(61*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(61*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[2*POS_CACHE_WIDTH-1:1*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(61*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(61*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[57*POS_CACHE_WIDTH-1:56*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(61*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(61*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[33*POS_CACHE_WIDTH-1:32*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(61*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(61*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[1*POS_CACHE_WIDTH-1:0*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(61*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(61*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[9*POS_CACHE_WIDTH-1:8*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(61*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(61*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[41*POS_CACHE_WIDTH-1:40*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(61*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(61*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[45*POS_CACHE_WIDTH-1:44*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(61*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(61*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[49*POS_CACHE_WIDTH-1:48*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(61*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(61*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[34*POS_CACHE_WIDTH-1:33*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(61*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(61*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[14*POS_CACHE_WIDTH-1:13*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(61*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(61*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[58*POS_CACHE_WIDTH-1:57*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(61*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(61*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[63*POS_CACHE_WIDTH-1:62*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(62*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(62*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[63*POS_CACHE_WIDTH-1:62*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(62*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(62*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[48*POS_CACHE_WIDTH-1:47*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(62*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(62*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[3*POS_CACHE_WIDTH-1:2*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(62*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(62*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[58*POS_CACHE_WIDTH-1:57*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(62*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(62*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[34*POS_CACHE_WIDTH-1:33*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(62*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(62*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[2*POS_CACHE_WIDTH-1:1*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(62*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(62*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[10*POS_CACHE_WIDTH-1:9*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(62*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(62*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[42*POS_CACHE_WIDTH-1:41*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(62*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(62*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[46*POS_CACHE_WIDTH-1:45*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(62*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(62*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[50*POS_CACHE_WIDTH-1:49*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(62*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(62*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[35*POS_CACHE_WIDTH-1:34*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(62*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(62*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[15*POS_CACHE_WIDTH-1:14*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(62*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(62*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[59*POS_CACHE_WIDTH-1:58*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(62*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(62*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[64*POS_CACHE_WIDTH-1:63*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(63*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH-1:(63*(NUM_NEIGHBOR_CELLS+1)+0)*POS_CACHE_WIDTH] = rd_nb_position[64*POS_CACHE_WIDTH-1:63*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(63*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH-1:(63*(NUM_NEIGHBOR_CELLS+1)+1)*POS_CACHE_WIDTH] = rd_nb_position[45*POS_CACHE_WIDTH-1:44*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(63*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH-1:(63*(NUM_NEIGHBOR_CELLS+1)+2)*POS_CACHE_WIDTH] = rd_nb_position[4*POS_CACHE_WIDTH-1:3*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(63*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH-1:(63*(NUM_NEIGHBOR_CELLS+1)+3)*POS_CACHE_WIDTH] = rd_nb_position[59*POS_CACHE_WIDTH-1:58*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(63*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH-1:(63*(NUM_NEIGHBOR_CELLS+1)+4)*POS_CACHE_WIDTH] = rd_nb_position[35*POS_CACHE_WIDTH-1:34*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(63*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH-1:(63*(NUM_NEIGHBOR_CELLS+1)+5)*POS_CACHE_WIDTH] = rd_nb_position[3*POS_CACHE_WIDTH-1:2*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(63*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH-1:(63*(NUM_NEIGHBOR_CELLS+1)+6)*POS_CACHE_WIDTH] = rd_nb_position[11*POS_CACHE_WIDTH-1:10*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(63*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH-1:(63*(NUM_NEIGHBOR_CELLS+1)+7)*POS_CACHE_WIDTH] = rd_nb_position[43*POS_CACHE_WIDTH-1:42*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(63*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH-1:(63*(NUM_NEIGHBOR_CELLS+1)+8)*POS_CACHE_WIDTH] = rd_nb_position[47*POS_CACHE_WIDTH-1:46*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(63*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH-1:(63*(NUM_NEIGHBOR_CELLS+1)+9)*POS_CACHE_WIDTH] = rd_nb_position[51*POS_CACHE_WIDTH-1:50*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(63*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH-1:(63*(NUM_NEIGHBOR_CELLS+1)+10)*POS_CACHE_WIDTH] = rd_nb_position[36*POS_CACHE_WIDTH-1:35*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(63*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH-1:(63*(NUM_NEIGHBOR_CELLS+1)+11)*POS_CACHE_WIDTH] = rd_nb_position[16*POS_CACHE_WIDTH-1:15*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(63*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH-1:(63*(NUM_NEIGHBOR_CELLS+1)+12)*POS_CACHE_WIDTH] = rd_nb_position[60*POS_CACHE_WIDTH-1:59*POS_CACHE_WIDTH];
assign rd_nb_position_splitted[(63*(NUM_NEIGHBOR_CELLS+1)+14)*POS_CACHE_WIDTH-1:(63*(NUM_NEIGHBOR_CELLS+1)+13)*POS_CACHE_WIDTH] = rd_nb_position[61*POS_CACHE_WIDTH-1:60*POS_CACHE_WIDTH];


assign broadcast_done_splitted[0*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[0];
assign broadcast_done_splitted[0*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[49];
assign broadcast_done_splitted[0*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[20];
assign broadcast_done_splitted[0*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[15];
assign broadcast_done_splitted[0*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[55];
assign broadcast_done_splitted[0*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[23];
assign broadcast_done_splitted[0*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[31];
assign broadcast_done_splitted[0*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[63];
assign broadcast_done_splitted[0*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[51];
assign broadcast_done_splitted[0*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[7];
assign broadcast_done_splitted[0*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[52];
assign broadcast_done_splitted[0*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[16];
assign broadcast_done_splitted[0*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[12];
assign broadcast_done_splitted[0*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[1];
assign broadcast_done_splitted[1*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[1];
assign broadcast_done_splitted[1*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[50];
assign broadcast_done_splitted[1*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[21];
assign broadcast_done_splitted[1*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[12];
assign broadcast_done_splitted[1*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[52];
assign broadcast_done_splitted[1*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[20];
assign broadcast_done_splitted[1*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[28];
assign broadcast_done_splitted[1*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[60];
assign broadcast_done_splitted[1*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[48];
assign broadcast_done_splitted[1*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[4];
assign broadcast_done_splitted[1*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[53];
assign broadcast_done_splitted[1*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[17];
assign broadcast_done_splitted[1*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[13];
assign broadcast_done_splitted[1*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[2];
assign broadcast_done_splitted[2*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[2];
assign broadcast_done_splitted[2*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[51];
assign broadcast_done_splitted[2*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[22];
assign broadcast_done_splitted[2*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[13];
assign broadcast_done_splitted[2*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[53];
assign broadcast_done_splitted[2*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[21];
assign broadcast_done_splitted[2*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[29];
assign broadcast_done_splitted[2*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[61];
assign broadcast_done_splitted[2*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[49];
assign broadcast_done_splitted[2*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[5];
assign broadcast_done_splitted[2*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[54];
assign broadcast_done_splitted[2*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[18];
assign broadcast_done_splitted[2*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[14];
assign broadcast_done_splitted[2*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[3];
assign broadcast_done_splitted[3*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[3];
assign broadcast_done_splitted[3*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[48];
assign broadcast_done_splitted[3*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[23];
assign broadcast_done_splitted[3*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[14];
assign broadcast_done_splitted[3*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[54];
assign broadcast_done_splitted[3*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[22];
assign broadcast_done_splitted[3*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[30];
assign broadcast_done_splitted[3*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[62];
assign broadcast_done_splitted[3*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[50];
assign broadcast_done_splitted[3*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[6];
assign broadcast_done_splitted[3*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[55];
assign broadcast_done_splitted[3*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[19];
assign broadcast_done_splitted[3*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[15];
assign broadcast_done_splitted[3*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[0];
assign broadcast_done_splitted[4*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[4];
assign broadcast_done_splitted[4*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[53];
assign broadcast_done_splitted[4*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[24];
assign broadcast_done_splitted[4*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[3];
assign broadcast_done_splitted[4*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[59];
assign broadcast_done_splitted[4*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[27];
assign broadcast_done_splitted[4*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[19];
assign broadcast_done_splitted[4*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[51];
assign broadcast_done_splitted[4*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[55];
assign broadcast_done_splitted[4*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[11];
assign broadcast_done_splitted[4*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[56];
assign broadcast_done_splitted[4*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[20];
assign broadcast_done_splitted[4*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[0];
assign broadcast_done_splitted[4*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[5];
assign broadcast_done_splitted[5*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[5];
assign broadcast_done_splitted[5*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[54];
assign broadcast_done_splitted[5*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[25];
assign broadcast_done_splitted[5*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[0];
assign broadcast_done_splitted[5*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[56];
assign broadcast_done_splitted[5*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[24];
assign broadcast_done_splitted[5*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[16];
assign broadcast_done_splitted[5*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[48];
assign broadcast_done_splitted[5*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[52];
assign broadcast_done_splitted[5*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[8];
assign broadcast_done_splitted[5*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[57];
assign broadcast_done_splitted[5*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[21];
assign broadcast_done_splitted[5*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[1];
assign broadcast_done_splitted[5*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[6];
assign broadcast_done_splitted[6*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[6];
assign broadcast_done_splitted[6*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[55];
assign broadcast_done_splitted[6*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[26];
assign broadcast_done_splitted[6*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[1];
assign broadcast_done_splitted[6*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[57];
assign broadcast_done_splitted[6*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[25];
assign broadcast_done_splitted[6*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[17];
assign broadcast_done_splitted[6*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[49];
assign broadcast_done_splitted[6*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[53];
assign broadcast_done_splitted[6*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[9];
assign broadcast_done_splitted[6*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[58];
assign broadcast_done_splitted[6*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[22];
assign broadcast_done_splitted[6*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[2];
assign broadcast_done_splitted[6*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[7];
assign broadcast_done_splitted[7*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[7];
assign broadcast_done_splitted[7*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[52];
assign broadcast_done_splitted[7*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[27];
assign broadcast_done_splitted[7*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[2];
assign broadcast_done_splitted[7*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[58];
assign broadcast_done_splitted[7*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[26];
assign broadcast_done_splitted[7*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[18];
assign broadcast_done_splitted[7*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[50];
assign broadcast_done_splitted[7*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[54];
assign broadcast_done_splitted[7*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[10];
assign broadcast_done_splitted[7*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[59];
assign broadcast_done_splitted[7*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[23];
assign broadcast_done_splitted[7*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[3];
assign broadcast_done_splitted[7*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[4];
assign broadcast_done_splitted[8*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[8];
assign broadcast_done_splitted[8*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[57];
assign broadcast_done_splitted[8*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[28];
assign broadcast_done_splitted[8*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[7];
assign broadcast_done_splitted[8*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[63];
assign broadcast_done_splitted[8*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[31];
assign broadcast_done_splitted[8*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[23];
assign broadcast_done_splitted[8*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[55];
assign broadcast_done_splitted[8*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[59];
assign broadcast_done_splitted[8*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[15];
assign broadcast_done_splitted[8*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[60];
assign broadcast_done_splitted[8*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[24];
assign broadcast_done_splitted[8*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[4];
assign broadcast_done_splitted[8*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[9];
assign broadcast_done_splitted[9*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[9];
assign broadcast_done_splitted[9*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[58];
assign broadcast_done_splitted[9*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[29];
assign broadcast_done_splitted[9*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[4];
assign broadcast_done_splitted[9*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[60];
assign broadcast_done_splitted[9*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[28];
assign broadcast_done_splitted[9*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[20];
assign broadcast_done_splitted[9*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[52];
assign broadcast_done_splitted[9*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[56];
assign broadcast_done_splitted[9*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[12];
assign broadcast_done_splitted[9*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[61];
assign broadcast_done_splitted[9*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[25];
assign broadcast_done_splitted[9*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[5];
assign broadcast_done_splitted[9*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[10];
assign broadcast_done_splitted[10*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[10];
assign broadcast_done_splitted[10*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[59];
assign broadcast_done_splitted[10*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[30];
assign broadcast_done_splitted[10*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[5];
assign broadcast_done_splitted[10*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[61];
assign broadcast_done_splitted[10*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[29];
assign broadcast_done_splitted[10*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[21];
assign broadcast_done_splitted[10*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[53];
assign broadcast_done_splitted[10*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[57];
assign broadcast_done_splitted[10*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[13];
assign broadcast_done_splitted[10*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[62];
assign broadcast_done_splitted[10*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[26];
assign broadcast_done_splitted[10*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[6];
assign broadcast_done_splitted[10*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[11];
assign broadcast_done_splitted[11*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[11];
assign broadcast_done_splitted[11*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[56];
assign broadcast_done_splitted[11*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[31];
assign broadcast_done_splitted[11*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[6];
assign broadcast_done_splitted[11*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[62];
assign broadcast_done_splitted[11*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[30];
assign broadcast_done_splitted[11*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[22];
assign broadcast_done_splitted[11*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[54];
assign broadcast_done_splitted[11*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[58];
assign broadcast_done_splitted[11*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[14];
assign broadcast_done_splitted[11*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[63];
assign broadcast_done_splitted[11*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[27];
assign broadcast_done_splitted[11*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[7];
assign broadcast_done_splitted[11*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[8];
assign broadcast_done_splitted[12*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[12];
assign broadcast_done_splitted[12*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[61];
assign broadcast_done_splitted[12*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[16];
assign broadcast_done_splitted[12*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[11];
assign broadcast_done_splitted[12*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[51];
assign broadcast_done_splitted[12*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[19];
assign broadcast_done_splitted[12*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[27];
assign broadcast_done_splitted[12*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[59];
assign broadcast_done_splitted[12*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[63];
assign broadcast_done_splitted[12*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[3];
assign broadcast_done_splitted[12*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[48];
assign broadcast_done_splitted[12*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[28];
assign broadcast_done_splitted[12*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[8];
assign broadcast_done_splitted[12*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[13];
assign broadcast_done_splitted[13*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[13];
assign broadcast_done_splitted[13*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[62];
assign broadcast_done_splitted[13*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[17];
assign broadcast_done_splitted[13*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[8];
assign broadcast_done_splitted[13*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[48];
assign broadcast_done_splitted[13*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[16];
assign broadcast_done_splitted[13*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[24];
assign broadcast_done_splitted[13*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[56];
assign broadcast_done_splitted[13*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[60];
assign broadcast_done_splitted[13*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[0];
assign broadcast_done_splitted[13*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[49];
assign broadcast_done_splitted[13*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[29];
assign broadcast_done_splitted[13*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[9];
assign broadcast_done_splitted[13*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[14];
assign broadcast_done_splitted[14*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[14];
assign broadcast_done_splitted[14*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[63];
assign broadcast_done_splitted[14*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[18];
assign broadcast_done_splitted[14*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[9];
assign broadcast_done_splitted[14*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[49];
assign broadcast_done_splitted[14*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[17];
assign broadcast_done_splitted[14*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[25];
assign broadcast_done_splitted[14*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[57];
assign broadcast_done_splitted[14*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[61];
assign broadcast_done_splitted[14*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[1];
assign broadcast_done_splitted[14*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[50];
assign broadcast_done_splitted[14*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[30];
assign broadcast_done_splitted[14*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[10];
assign broadcast_done_splitted[14*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[15];
assign broadcast_done_splitted[15*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[15];
assign broadcast_done_splitted[15*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[60];
assign broadcast_done_splitted[15*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[19];
assign broadcast_done_splitted[15*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[10];
assign broadcast_done_splitted[15*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[50];
assign broadcast_done_splitted[15*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[18];
assign broadcast_done_splitted[15*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[26];
assign broadcast_done_splitted[15*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[58];
assign broadcast_done_splitted[15*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[62];
assign broadcast_done_splitted[15*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[2];
assign broadcast_done_splitted[15*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[51];
assign broadcast_done_splitted[15*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[31];
assign broadcast_done_splitted[15*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[11];
assign broadcast_done_splitted[15*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[12];
assign broadcast_done_splitted[16*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[16];
assign broadcast_done_splitted[16*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[1];
assign broadcast_done_splitted[16*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[36];
assign broadcast_done_splitted[16*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[31];
assign broadcast_done_splitted[16*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[7];
assign broadcast_done_splitted[16*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[39];
assign broadcast_done_splitted[16*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[47];
assign broadcast_done_splitted[16*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[15];
assign broadcast_done_splitted[16*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[3];
assign broadcast_done_splitted[16*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[23];
assign broadcast_done_splitted[16*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[4];
assign broadcast_done_splitted[16*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[32];
assign broadcast_done_splitted[16*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[28];
assign broadcast_done_splitted[16*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[17];
assign broadcast_done_splitted[17*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[17];
assign broadcast_done_splitted[17*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[2];
assign broadcast_done_splitted[17*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[37];
assign broadcast_done_splitted[17*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[28];
assign broadcast_done_splitted[17*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[4];
assign broadcast_done_splitted[17*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[36];
assign broadcast_done_splitted[17*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[44];
assign broadcast_done_splitted[17*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[12];
assign broadcast_done_splitted[17*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[0];
assign broadcast_done_splitted[17*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[20];
assign broadcast_done_splitted[17*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[5];
assign broadcast_done_splitted[17*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[33];
assign broadcast_done_splitted[17*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[29];
assign broadcast_done_splitted[17*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[18];
assign broadcast_done_splitted[18*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[18];
assign broadcast_done_splitted[18*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[3];
assign broadcast_done_splitted[18*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[38];
assign broadcast_done_splitted[18*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[29];
assign broadcast_done_splitted[18*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[5];
assign broadcast_done_splitted[18*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[37];
assign broadcast_done_splitted[18*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[45];
assign broadcast_done_splitted[18*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[13];
assign broadcast_done_splitted[18*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[1];
assign broadcast_done_splitted[18*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[21];
assign broadcast_done_splitted[18*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[6];
assign broadcast_done_splitted[18*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[34];
assign broadcast_done_splitted[18*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[30];
assign broadcast_done_splitted[18*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[19];
assign broadcast_done_splitted[19*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[19];
assign broadcast_done_splitted[19*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[0];
assign broadcast_done_splitted[19*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[39];
assign broadcast_done_splitted[19*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[30];
assign broadcast_done_splitted[19*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[6];
assign broadcast_done_splitted[19*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[38];
assign broadcast_done_splitted[19*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[46];
assign broadcast_done_splitted[19*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[14];
assign broadcast_done_splitted[19*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[2];
assign broadcast_done_splitted[19*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[22];
assign broadcast_done_splitted[19*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[7];
assign broadcast_done_splitted[19*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[35];
assign broadcast_done_splitted[19*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[31];
assign broadcast_done_splitted[19*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[16];
assign broadcast_done_splitted[20*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[20];
assign broadcast_done_splitted[20*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[5];
assign broadcast_done_splitted[20*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[40];
assign broadcast_done_splitted[20*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[19];
assign broadcast_done_splitted[20*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[11];
assign broadcast_done_splitted[20*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[43];
assign broadcast_done_splitted[20*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[35];
assign broadcast_done_splitted[20*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[3];
assign broadcast_done_splitted[20*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[7];
assign broadcast_done_splitted[20*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[27];
assign broadcast_done_splitted[20*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[8];
assign broadcast_done_splitted[20*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[36];
assign broadcast_done_splitted[20*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[16];
assign broadcast_done_splitted[20*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[21];
assign broadcast_done_splitted[21*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[21];
assign broadcast_done_splitted[21*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[6];
assign broadcast_done_splitted[21*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[41];
assign broadcast_done_splitted[21*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[16];
assign broadcast_done_splitted[21*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[8];
assign broadcast_done_splitted[21*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[40];
assign broadcast_done_splitted[21*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[32];
assign broadcast_done_splitted[21*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[0];
assign broadcast_done_splitted[21*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[4];
assign broadcast_done_splitted[21*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[24];
assign broadcast_done_splitted[21*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[9];
assign broadcast_done_splitted[21*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[37];
assign broadcast_done_splitted[21*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[17];
assign broadcast_done_splitted[21*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[22];
assign broadcast_done_splitted[22*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[22];
assign broadcast_done_splitted[22*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[7];
assign broadcast_done_splitted[22*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[42];
assign broadcast_done_splitted[22*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[17];
assign broadcast_done_splitted[22*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[9];
assign broadcast_done_splitted[22*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[41];
assign broadcast_done_splitted[22*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[33];
assign broadcast_done_splitted[22*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[1];
assign broadcast_done_splitted[22*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[5];
assign broadcast_done_splitted[22*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[25];
assign broadcast_done_splitted[22*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[10];
assign broadcast_done_splitted[22*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[38];
assign broadcast_done_splitted[22*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[18];
assign broadcast_done_splitted[22*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[23];
assign broadcast_done_splitted[23*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[23];
assign broadcast_done_splitted[23*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[4];
assign broadcast_done_splitted[23*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[43];
assign broadcast_done_splitted[23*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[18];
assign broadcast_done_splitted[23*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[10];
assign broadcast_done_splitted[23*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[42];
assign broadcast_done_splitted[23*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[34];
assign broadcast_done_splitted[23*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[2];
assign broadcast_done_splitted[23*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[6];
assign broadcast_done_splitted[23*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[26];
assign broadcast_done_splitted[23*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[11];
assign broadcast_done_splitted[23*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[39];
assign broadcast_done_splitted[23*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[19];
assign broadcast_done_splitted[23*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[20];
assign broadcast_done_splitted[24*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[24];
assign broadcast_done_splitted[24*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[9];
assign broadcast_done_splitted[24*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[44];
assign broadcast_done_splitted[24*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[23];
assign broadcast_done_splitted[24*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[15];
assign broadcast_done_splitted[24*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[47];
assign broadcast_done_splitted[24*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[39];
assign broadcast_done_splitted[24*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[7];
assign broadcast_done_splitted[24*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[11];
assign broadcast_done_splitted[24*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[31];
assign broadcast_done_splitted[24*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[12];
assign broadcast_done_splitted[24*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[40];
assign broadcast_done_splitted[24*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[20];
assign broadcast_done_splitted[24*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[25];
assign broadcast_done_splitted[25*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[25];
assign broadcast_done_splitted[25*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[10];
assign broadcast_done_splitted[25*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[45];
assign broadcast_done_splitted[25*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[20];
assign broadcast_done_splitted[25*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[12];
assign broadcast_done_splitted[25*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[44];
assign broadcast_done_splitted[25*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[36];
assign broadcast_done_splitted[25*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[4];
assign broadcast_done_splitted[25*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[8];
assign broadcast_done_splitted[25*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[28];
assign broadcast_done_splitted[25*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[13];
assign broadcast_done_splitted[25*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[41];
assign broadcast_done_splitted[25*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[21];
assign broadcast_done_splitted[25*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[26];
assign broadcast_done_splitted[26*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[26];
assign broadcast_done_splitted[26*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[11];
assign broadcast_done_splitted[26*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[46];
assign broadcast_done_splitted[26*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[21];
assign broadcast_done_splitted[26*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[13];
assign broadcast_done_splitted[26*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[45];
assign broadcast_done_splitted[26*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[37];
assign broadcast_done_splitted[26*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[5];
assign broadcast_done_splitted[26*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[9];
assign broadcast_done_splitted[26*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[29];
assign broadcast_done_splitted[26*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[14];
assign broadcast_done_splitted[26*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[42];
assign broadcast_done_splitted[26*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[22];
assign broadcast_done_splitted[26*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[27];
assign broadcast_done_splitted[27*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[27];
assign broadcast_done_splitted[27*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[8];
assign broadcast_done_splitted[27*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[47];
assign broadcast_done_splitted[27*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[22];
assign broadcast_done_splitted[27*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[14];
assign broadcast_done_splitted[27*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[46];
assign broadcast_done_splitted[27*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[38];
assign broadcast_done_splitted[27*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[6];
assign broadcast_done_splitted[27*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[10];
assign broadcast_done_splitted[27*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[30];
assign broadcast_done_splitted[27*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[15];
assign broadcast_done_splitted[27*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[43];
assign broadcast_done_splitted[27*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[23];
assign broadcast_done_splitted[27*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[24];
assign broadcast_done_splitted[28*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[28];
assign broadcast_done_splitted[28*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[13];
assign broadcast_done_splitted[28*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[32];
assign broadcast_done_splitted[28*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[27];
assign broadcast_done_splitted[28*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[3];
assign broadcast_done_splitted[28*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[35];
assign broadcast_done_splitted[28*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[43];
assign broadcast_done_splitted[28*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[11];
assign broadcast_done_splitted[28*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[15];
assign broadcast_done_splitted[28*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[19];
assign broadcast_done_splitted[28*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[0];
assign broadcast_done_splitted[28*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[44];
assign broadcast_done_splitted[28*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[24];
assign broadcast_done_splitted[28*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[29];
assign broadcast_done_splitted[29*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[29];
assign broadcast_done_splitted[29*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[14];
assign broadcast_done_splitted[29*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[33];
assign broadcast_done_splitted[29*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[24];
assign broadcast_done_splitted[29*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[0];
assign broadcast_done_splitted[29*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[32];
assign broadcast_done_splitted[29*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[40];
assign broadcast_done_splitted[29*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[8];
assign broadcast_done_splitted[29*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[12];
assign broadcast_done_splitted[29*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[16];
assign broadcast_done_splitted[29*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[1];
assign broadcast_done_splitted[29*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[45];
assign broadcast_done_splitted[29*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[25];
assign broadcast_done_splitted[29*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[30];
assign broadcast_done_splitted[30*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[30];
assign broadcast_done_splitted[30*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[15];
assign broadcast_done_splitted[30*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[34];
assign broadcast_done_splitted[30*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[25];
assign broadcast_done_splitted[30*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[1];
assign broadcast_done_splitted[30*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[33];
assign broadcast_done_splitted[30*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[41];
assign broadcast_done_splitted[30*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[9];
assign broadcast_done_splitted[30*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[13];
assign broadcast_done_splitted[30*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[17];
assign broadcast_done_splitted[30*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[2];
assign broadcast_done_splitted[30*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[46];
assign broadcast_done_splitted[30*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[26];
assign broadcast_done_splitted[30*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[31];
assign broadcast_done_splitted[31*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[31];
assign broadcast_done_splitted[31*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[12];
assign broadcast_done_splitted[31*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[35];
assign broadcast_done_splitted[31*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[26];
assign broadcast_done_splitted[31*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[2];
assign broadcast_done_splitted[31*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[34];
assign broadcast_done_splitted[31*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[42];
assign broadcast_done_splitted[31*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[10];
assign broadcast_done_splitted[31*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[14];
assign broadcast_done_splitted[31*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[18];
assign broadcast_done_splitted[31*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[3];
assign broadcast_done_splitted[31*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[47];
assign broadcast_done_splitted[31*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[27];
assign broadcast_done_splitted[31*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[28];
assign broadcast_done_splitted[32*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[32];
assign broadcast_done_splitted[32*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[17];
assign broadcast_done_splitted[32*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[52];
assign broadcast_done_splitted[32*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[47];
assign broadcast_done_splitted[32*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[23];
assign broadcast_done_splitted[32*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[55];
assign broadcast_done_splitted[32*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[63];
assign broadcast_done_splitted[32*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[31];
assign broadcast_done_splitted[32*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[19];
assign broadcast_done_splitted[32*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[39];
assign broadcast_done_splitted[32*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[20];
assign broadcast_done_splitted[32*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[48];
assign broadcast_done_splitted[32*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[44];
assign broadcast_done_splitted[32*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[33];
assign broadcast_done_splitted[33*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[33];
assign broadcast_done_splitted[33*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[18];
assign broadcast_done_splitted[33*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[53];
assign broadcast_done_splitted[33*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[44];
assign broadcast_done_splitted[33*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[20];
assign broadcast_done_splitted[33*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[52];
assign broadcast_done_splitted[33*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[60];
assign broadcast_done_splitted[33*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[28];
assign broadcast_done_splitted[33*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[16];
assign broadcast_done_splitted[33*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[36];
assign broadcast_done_splitted[33*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[21];
assign broadcast_done_splitted[33*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[49];
assign broadcast_done_splitted[33*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[45];
assign broadcast_done_splitted[33*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[34];
assign broadcast_done_splitted[34*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[34];
assign broadcast_done_splitted[34*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[19];
assign broadcast_done_splitted[34*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[54];
assign broadcast_done_splitted[34*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[45];
assign broadcast_done_splitted[34*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[21];
assign broadcast_done_splitted[34*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[53];
assign broadcast_done_splitted[34*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[61];
assign broadcast_done_splitted[34*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[29];
assign broadcast_done_splitted[34*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[17];
assign broadcast_done_splitted[34*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[37];
assign broadcast_done_splitted[34*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[22];
assign broadcast_done_splitted[34*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[50];
assign broadcast_done_splitted[34*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[46];
assign broadcast_done_splitted[34*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[35];
assign broadcast_done_splitted[35*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[35];
assign broadcast_done_splitted[35*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[16];
assign broadcast_done_splitted[35*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[55];
assign broadcast_done_splitted[35*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[46];
assign broadcast_done_splitted[35*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[22];
assign broadcast_done_splitted[35*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[54];
assign broadcast_done_splitted[35*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[62];
assign broadcast_done_splitted[35*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[30];
assign broadcast_done_splitted[35*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[18];
assign broadcast_done_splitted[35*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[38];
assign broadcast_done_splitted[35*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[23];
assign broadcast_done_splitted[35*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[51];
assign broadcast_done_splitted[35*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[47];
assign broadcast_done_splitted[35*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[32];
assign broadcast_done_splitted[36*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[36];
assign broadcast_done_splitted[36*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[21];
assign broadcast_done_splitted[36*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[56];
assign broadcast_done_splitted[36*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[35];
assign broadcast_done_splitted[36*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[27];
assign broadcast_done_splitted[36*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[59];
assign broadcast_done_splitted[36*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[51];
assign broadcast_done_splitted[36*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[19];
assign broadcast_done_splitted[36*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[23];
assign broadcast_done_splitted[36*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[43];
assign broadcast_done_splitted[36*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[24];
assign broadcast_done_splitted[36*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[52];
assign broadcast_done_splitted[36*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[32];
assign broadcast_done_splitted[36*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[37];
assign broadcast_done_splitted[37*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[37];
assign broadcast_done_splitted[37*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[22];
assign broadcast_done_splitted[37*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[57];
assign broadcast_done_splitted[37*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[32];
assign broadcast_done_splitted[37*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[24];
assign broadcast_done_splitted[37*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[56];
assign broadcast_done_splitted[37*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[48];
assign broadcast_done_splitted[37*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[16];
assign broadcast_done_splitted[37*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[20];
assign broadcast_done_splitted[37*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[40];
assign broadcast_done_splitted[37*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[25];
assign broadcast_done_splitted[37*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[53];
assign broadcast_done_splitted[37*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[33];
assign broadcast_done_splitted[37*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[38];
assign broadcast_done_splitted[38*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[38];
assign broadcast_done_splitted[38*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[23];
assign broadcast_done_splitted[38*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[58];
assign broadcast_done_splitted[38*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[33];
assign broadcast_done_splitted[38*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[25];
assign broadcast_done_splitted[38*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[57];
assign broadcast_done_splitted[38*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[49];
assign broadcast_done_splitted[38*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[17];
assign broadcast_done_splitted[38*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[21];
assign broadcast_done_splitted[38*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[41];
assign broadcast_done_splitted[38*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[26];
assign broadcast_done_splitted[38*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[54];
assign broadcast_done_splitted[38*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[34];
assign broadcast_done_splitted[38*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[39];
assign broadcast_done_splitted[39*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[39];
assign broadcast_done_splitted[39*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[20];
assign broadcast_done_splitted[39*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[59];
assign broadcast_done_splitted[39*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[34];
assign broadcast_done_splitted[39*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[26];
assign broadcast_done_splitted[39*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[58];
assign broadcast_done_splitted[39*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[50];
assign broadcast_done_splitted[39*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[18];
assign broadcast_done_splitted[39*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[22];
assign broadcast_done_splitted[39*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[42];
assign broadcast_done_splitted[39*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[27];
assign broadcast_done_splitted[39*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[55];
assign broadcast_done_splitted[39*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[35];
assign broadcast_done_splitted[39*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[36];
assign broadcast_done_splitted[40*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[40];
assign broadcast_done_splitted[40*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[25];
assign broadcast_done_splitted[40*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[60];
assign broadcast_done_splitted[40*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[39];
assign broadcast_done_splitted[40*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[31];
assign broadcast_done_splitted[40*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[63];
assign broadcast_done_splitted[40*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[55];
assign broadcast_done_splitted[40*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[23];
assign broadcast_done_splitted[40*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[27];
assign broadcast_done_splitted[40*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[47];
assign broadcast_done_splitted[40*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[28];
assign broadcast_done_splitted[40*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[56];
assign broadcast_done_splitted[40*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[36];
assign broadcast_done_splitted[40*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[41];
assign broadcast_done_splitted[41*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[41];
assign broadcast_done_splitted[41*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[26];
assign broadcast_done_splitted[41*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[61];
assign broadcast_done_splitted[41*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[36];
assign broadcast_done_splitted[41*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[28];
assign broadcast_done_splitted[41*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[60];
assign broadcast_done_splitted[41*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[52];
assign broadcast_done_splitted[41*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[20];
assign broadcast_done_splitted[41*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[24];
assign broadcast_done_splitted[41*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[44];
assign broadcast_done_splitted[41*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[29];
assign broadcast_done_splitted[41*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[57];
assign broadcast_done_splitted[41*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[37];
assign broadcast_done_splitted[41*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[42];
assign broadcast_done_splitted[42*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[42];
assign broadcast_done_splitted[42*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[27];
assign broadcast_done_splitted[42*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[62];
assign broadcast_done_splitted[42*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[37];
assign broadcast_done_splitted[42*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[29];
assign broadcast_done_splitted[42*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[61];
assign broadcast_done_splitted[42*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[53];
assign broadcast_done_splitted[42*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[21];
assign broadcast_done_splitted[42*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[25];
assign broadcast_done_splitted[42*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[45];
assign broadcast_done_splitted[42*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[30];
assign broadcast_done_splitted[42*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[58];
assign broadcast_done_splitted[42*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[38];
assign broadcast_done_splitted[42*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[43];
assign broadcast_done_splitted[43*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[43];
assign broadcast_done_splitted[43*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[24];
assign broadcast_done_splitted[43*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[63];
assign broadcast_done_splitted[43*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[38];
assign broadcast_done_splitted[43*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[30];
assign broadcast_done_splitted[43*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[62];
assign broadcast_done_splitted[43*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[54];
assign broadcast_done_splitted[43*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[22];
assign broadcast_done_splitted[43*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[26];
assign broadcast_done_splitted[43*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[46];
assign broadcast_done_splitted[43*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[31];
assign broadcast_done_splitted[43*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[59];
assign broadcast_done_splitted[43*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[39];
assign broadcast_done_splitted[43*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[40];
assign broadcast_done_splitted[44*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[44];
assign broadcast_done_splitted[44*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[29];
assign broadcast_done_splitted[44*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[48];
assign broadcast_done_splitted[44*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[43];
assign broadcast_done_splitted[44*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[19];
assign broadcast_done_splitted[44*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[51];
assign broadcast_done_splitted[44*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[59];
assign broadcast_done_splitted[44*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[27];
assign broadcast_done_splitted[44*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[31];
assign broadcast_done_splitted[44*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[35];
assign broadcast_done_splitted[44*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[16];
assign broadcast_done_splitted[44*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[60];
assign broadcast_done_splitted[44*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[40];
assign broadcast_done_splitted[44*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[45];
assign broadcast_done_splitted[45*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[45];
assign broadcast_done_splitted[45*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[30];
assign broadcast_done_splitted[45*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[49];
assign broadcast_done_splitted[45*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[40];
assign broadcast_done_splitted[45*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[16];
assign broadcast_done_splitted[45*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[48];
assign broadcast_done_splitted[45*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[56];
assign broadcast_done_splitted[45*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[24];
assign broadcast_done_splitted[45*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[28];
assign broadcast_done_splitted[45*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[32];
assign broadcast_done_splitted[45*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[17];
assign broadcast_done_splitted[45*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[61];
assign broadcast_done_splitted[45*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[41];
assign broadcast_done_splitted[45*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[46];
assign broadcast_done_splitted[46*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[46];
assign broadcast_done_splitted[46*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[31];
assign broadcast_done_splitted[46*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[50];
assign broadcast_done_splitted[46*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[41];
assign broadcast_done_splitted[46*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[17];
assign broadcast_done_splitted[46*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[49];
assign broadcast_done_splitted[46*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[57];
assign broadcast_done_splitted[46*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[25];
assign broadcast_done_splitted[46*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[29];
assign broadcast_done_splitted[46*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[33];
assign broadcast_done_splitted[46*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[18];
assign broadcast_done_splitted[46*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[62];
assign broadcast_done_splitted[46*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[42];
assign broadcast_done_splitted[46*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[47];
assign broadcast_done_splitted[47*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[47];
assign broadcast_done_splitted[47*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[28];
assign broadcast_done_splitted[47*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[51];
assign broadcast_done_splitted[47*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[42];
assign broadcast_done_splitted[47*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[18];
assign broadcast_done_splitted[47*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[50];
assign broadcast_done_splitted[47*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[58];
assign broadcast_done_splitted[47*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[26];
assign broadcast_done_splitted[47*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[30];
assign broadcast_done_splitted[47*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[34];
assign broadcast_done_splitted[47*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[19];
assign broadcast_done_splitted[47*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[63];
assign broadcast_done_splitted[47*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[43];
assign broadcast_done_splitted[47*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[44];
assign broadcast_done_splitted[48*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[48];
assign broadcast_done_splitted[48*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[33];
assign broadcast_done_splitted[48*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[4];
assign broadcast_done_splitted[48*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[63];
assign broadcast_done_splitted[48*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[39];
assign broadcast_done_splitted[48*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[7];
assign broadcast_done_splitted[48*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[15];
assign broadcast_done_splitted[48*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[47];
assign broadcast_done_splitted[48*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[35];
assign broadcast_done_splitted[48*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[55];
assign broadcast_done_splitted[48*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[36];
assign broadcast_done_splitted[48*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[0];
assign broadcast_done_splitted[48*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[60];
assign broadcast_done_splitted[48*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[49];
assign broadcast_done_splitted[49*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[49];
assign broadcast_done_splitted[49*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[34];
assign broadcast_done_splitted[49*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[5];
assign broadcast_done_splitted[49*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[60];
assign broadcast_done_splitted[49*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[36];
assign broadcast_done_splitted[49*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[4];
assign broadcast_done_splitted[49*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[12];
assign broadcast_done_splitted[49*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[44];
assign broadcast_done_splitted[49*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[32];
assign broadcast_done_splitted[49*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[52];
assign broadcast_done_splitted[49*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[37];
assign broadcast_done_splitted[49*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[1];
assign broadcast_done_splitted[49*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[61];
assign broadcast_done_splitted[49*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[50];
assign broadcast_done_splitted[50*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[50];
assign broadcast_done_splitted[50*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[35];
assign broadcast_done_splitted[50*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[6];
assign broadcast_done_splitted[50*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[61];
assign broadcast_done_splitted[50*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[37];
assign broadcast_done_splitted[50*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[5];
assign broadcast_done_splitted[50*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[13];
assign broadcast_done_splitted[50*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[45];
assign broadcast_done_splitted[50*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[33];
assign broadcast_done_splitted[50*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[53];
assign broadcast_done_splitted[50*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[38];
assign broadcast_done_splitted[50*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[2];
assign broadcast_done_splitted[50*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[62];
assign broadcast_done_splitted[50*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[51];
assign broadcast_done_splitted[51*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[51];
assign broadcast_done_splitted[51*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[32];
assign broadcast_done_splitted[51*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[7];
assign broadcast_done_splitted[51*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[62];
assign broadcast_done_splitted[51*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[38];
assign broadcast_done_splitted[51*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[6];
assign broadcast_done_splitted[51*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[14];
assign broadcast_done_splitted[51*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[46];
assign broadcast_done_splitted[51*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[34];
assign broadcast_done_splitted[51*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[54];
assign broadcast_done_splitted[51*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[39];
assign broadcast_done_splitted[51*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[3];
assign broadcast_done_splitted[51*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[63];
assign broadcast_done_splitted[51*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[48];
assign broadcast_done_splitted[52*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[52];
assign broadcast_done_splitted[52*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[37];
assign broadcast_done_splitted[52*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[8];
assign broadcast_done_splitted[52*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[51];
assign broadcast_done_splitted[52*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[43];
assign broadcast_done_splitted[52*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[11];
assign broadcast_done_splitted[52*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[3];
assign broadcast_done_splitted[52*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[35];
assign broadcast_done_splitted[52*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[39];
assign broadcast_done_splitted[52*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[59];
assign broadcast_done_splitted[52*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[40];
assign broadcast_done_splitted[52*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[4];
assign broadcast_done_splitted[52*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[48];
assign broadcast_done_splitted[52*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[53];
assign broadcast_done_splitted[53*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[53];
assign broadcast_done_splitted[53*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[38];
assign broadcast_done_splitted[53*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[9];
assign broadcast_done_splitted[53*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[48];
assign broadcast_done_splitted[53*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[40];
assign broadcast_done_splitted[53*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[8];
assign broadcast_done_splitted[53*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[0];
assign broadcast_done_splitted[53*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[32];
assign broadcast_done_splitted[53*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[36];
assign broadcast_done_splitted[53*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[56];
assign broadcast_done_splitted[53*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[41];
assign broadcast_done_splitted[53*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[5];
assign broadcast_done_splitted[53*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[49];
assign broadcast_done_splitted[53*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[54];
assign broadcast_done_splitted[54*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[54];
assign broadcast_done_splitted[54*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[39];
assign broadcast_done_splitted[54*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[10];
assign broadcast_done_splitted[54*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[49];
assign broadcast_done_splitted[54*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[41];
assign broadcast_done_splitted[54*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[9];
assign broadcast_done_splitted[54*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[1];
assign broadcast_done_splitted[54*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[33];
assign broadcast_done_splitted[54*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[37];
assign broadcast_done_splitted[54*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[57];
assign broadcast_done_splitted[54*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[42];
assign broadcast_done_splitted[54*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[6];
assign broadcast_done_splitted[54*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[50];
assign broadcast_done_splitted[54*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[55];
assign broadcast_done_splitted[55*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[55];
assign broadcast_done_splitted[55*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[36];
assign broadcast_done_splitted[55*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[11];
assign broadcast_done_splitted[55*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[50];
assign broadcast_done_splitted[55*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[42];
assign broadcast_done_splitted[55*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[10];
assign broadcast_done_splitted[55*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[2];
assign broadcast_done_splitted[55*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[34];
assign broadcast_done_splitted[55*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[38];
assign broadcast_done_splitted[55*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[58];
assign broadcast_done_splitted[55*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[43];
assign broadcast_done_splitted[55*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[7];
assign broadcast_done_splitted[55*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[51];
assign broadcast_done_splitted[55*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[52];
assign broadcast_done_splitted[56*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[56];
assign broadcast_done_splitted[56*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[41];
assign broadcast_done_splitted[56*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[12];
assign broadcast_done_splitted[56*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[55];
assign broadcast_done_splitted[56*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[47];
assign broadcast_done_splitted[56*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[15];
assign broadcast_done_splitted[56*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[7];
assign broadcast_done_splitted[56*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[39];
assign broadcast_done_splitted[56*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[43];
assign broadcast_done_splitted[56*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[63];
assign broadcast_done_splitted[56*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[44];
assign broadcast_done_splitted[56*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[8];
assign broadcast_done_splitted[56*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[52];
assign broadcast_done_splitted[56*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[57];
assign broadcast_done_splitted[57*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[57];
assign broadcast_done_splitted[57*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[42];
assign broadcast_done_splitted[57*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[13];
assign broadcast_done_splitted[57*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[52];
assign broadcast_done_splitted[57*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[44];
assign broadcast_done_splitted[57*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[12];
assign broadcast_done_splitted[57*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[4];
assign broadcast_done_splitted[57*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[36];
assign broadcast_done_splitted[57*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[40];
assign broadcast_done_splitted[57*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[60];
assign broadcast_done_splitted[57*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[45];
assign broadcast_done_splitted[57*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[9];
assign broadcast_done_splitted[57*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[53];
assign broadcast_done_splitted[57*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[58];
assign broadcast_done_splitted[58*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[58];
assign broadcast_done_splitted[58*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[43];
assign broadcast_done_splitted[58*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[14];
assign broadcast_done_splitted[58*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[53];
assign broadcast_done_splitted[58*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[45];
assign broadcast_done_splitted[58*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[13];
assign broadcast_done_splitted[58*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[5];
assign broadcast_done_splitted[58*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[37];
assign broadcast_done_splitted[58*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[41];
assign broadcast_done_splitted[58*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[61];
assign broadcast_done_splitted[58*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[46];
assign broadcast_done_splitted[58*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[10];
assign broadcast_done_splitted[58*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[54];
assign broadcast_done_splitted[58*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[59];
assign broadcast_done_splitted[59*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[59];
assign broadcast_done_splitted[59*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[40];
assign broadcast_done_splitted[59*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[15];
assign broadcast_done_splitted[59*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[54];
assign broadcast_done_splitted[59*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[46];
assign broadcast_done_splitted[59*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[14];
assign broadcast_done_splitted[59*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[6];
assign broadcast_done_splitted[59*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[38];
assign broadcast_done_splitted[59*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[42];
assign broadcast_done_splitted[59*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[62];
assign broadcast_done_splitted[59*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[47];
assign broadcast_done_splitted[59*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[11];
assign broadcast_done_splitted[59*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[55];
assign broadcast_done_splitted[59*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[56];
assign broadcast_done_splitted[60*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[60];
assign broadcast_done_splitted[60*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[45];
assign broadcast_done_splitted[60*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[0];
assign broadcast_done_splitted[60*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[59];
assign broadcast_done_splitted[60*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[35];
assign broadcast_done_splitted[60*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[3];
assign broadcast_done_splitted[60*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[11];
assign broadcast_done_splitted[60*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[43];
assign broadcast_done_splitted[60*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[47];
assign broadcast_done_splitted[60*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[51];
assign broadcast_done_splitted[60*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[32];
assign broadcast_done_splitted[60*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[12];
assign broadcast_done_splitted[60*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[56];
assign broadcast_done_splitted[60*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[61];
assign broadcast_done_splitted[61*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[61];
assign broadcast_done_splitted[61*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[46];
assign broadcast_done_splitted[61*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[1];
assign broadcast_done_splitted[61*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[56];
assign broadcast_done_splitted[61*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[32];
assign broadcast_done_splitted[61*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[0];
assign broadcast_done_splitted[61*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[8];
assign broadcast_done_splitted[61*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[40];
assign broadcast_done_splitted[61*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[44];
assign broadcast_done_splitted[61*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[48];
assign broadcast_done_splitted[61*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[33];
assign broadcast_done_splitted[61*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[13];
assign broadcast_done_splitted[61*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[57];
assign broadcast_done_splitted[61*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[62];
assign broadcast_done_splitted[62*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[62];
assign broadcast_done_splitted[62*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[47];
assign broadcast_done_splitted[62*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[2];
assign broadcast_done_splitted[62*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[57];
assign broadcast_done_splitted[62*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[33];
assign broadcast_done_splitted[62*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[1];
assign broadcast_done_splitted[62*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[9];
assign broadcast_done_splitted[62*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[41];
assign broadcast_done_splitted[62*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[45];
assign broadcast_done_splitted[62*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[49];
assign broadcast_done_splitted[62*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[34];
assign broadcast_done_splitted[62*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[14];
assign broadcast_done_splitted[62*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[58];
assign broadcast_done_splitted[62*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[63];
assign broadcast_done_splitted[63*(NUM_NEIGHBOR_CELLS+1)+0] = broadcast_done[63];
assign broadcast_done_splitted[63*(NUM_NEIGHBOR_CELLS+1)+1] = broadcast_done[44];
assign broadcast_done_splitted[63*(NUM_NEIGHBOR_CELLS+1)+2] = broadcast_done[3];
assign broadcast_done_splitted[63*(NUM_NEIGHBOR_CELLS+1)+3] = broadcast_done[58];
assign broadcast_done_splitted[63*(NUM_NEIGHBOR_CELLS+1)+4] = broadcast_done[34];
assign broadcast_done_splitted[63*(NUM_NEIGHBOR_CELLS+1)+5] = broadcast_done[2];
assign broadcast_done_splitted[63*(NUM_NEIGHBOR_CELLS+1)+6] = broadcast_done[10];
assign broadcast_done_splitted[63*(NUM_NEIGHBOR_CELLS+1)+7] = broadcast_done[42];
assign broadcast_done_splitted[63*(NUM_NEIGHBOR_CELLS+1)+8] = broadcast_done[46];
assign broadcast_done_splitted[63*(NUM_NEIGHBOR_CELLS+1)+9] = broadcast_done[50];
assign broadcast_done_splitted[63*(NUM_NEIGHBOR_CELLS+1)+10] = broadcast_done[35];
assign broadcast_done_splitted[63*(NUM_NEIGHBOR_CELLS+1)+11] = broadcast_done[15];
assign broadcast_done_splitted[63*(NUM_NEIGHBOR_CELLS+1)+12] = broadcast_done[59];
assign broadcast_done_splitted[63*(NUM_NEIGHBOR_CELLS+1)+13] = broadcast_done[60];

endmodule