module single_cell_reading_pos_caches
#(
	parameter OFFSET_WIDTH = 29,
	parameter DATA_WIDTH = 3*OFFSET_WIDTH, 
	parameter PARTICLE_NUM = 127,
	parameter NUM_NEIGHBOR_CELLS = 13, 
	parameter ADDR_WIDTH = 7
)
(
	input clk,
	input [ADDR_WIDTH-1:0] particle_id, 
	output [(NUM_NEIGHBOR_CELLS+1)*DATA_WIDTH-1:0] pos_data
);

cell_2_2_2
#(
	.DATA_WIDTH(DATA_WIDTH), 
	.PARTICLE_NUM(PARTICLE_NUM), 
	.ADDR_WIDTH(7)
)
pos_cache_2_2_2
(
	.address(particle_id), 
	.clock(clk), 
	.data(), 
	.rden(1'b1), 
	.wren(1'b0), 
	.q(pos_data[DATA_WIDTH-1:0])
);
cell_2_2_3
#(
	.DATA_WIDTH(DATA_WIDTH), 
	.PARTICLE_NUM(PARTICLE_NUM), 
	.ADDR_WIDTH(7)
)
pos_cache_2_2_3
(
	.address(particle_id), 
	.clock(clk), 
	.data(), 
	.rden(1'b1), 
	.wren(1'b0), 
	.q(pos_data[2*DATA_WIDTH-1:DATA_WIDTH])
);
cell_2_3_1
#(
	.DATA_WIDTH(DATA_WIDTH), 
	.PARTICLE_NUM(PARTICLE_NUM), 
	.ADDR_WIDTH(7)
)
pos_cache_2_3_1
(
	.address(particle_id), 
	.clock(clk), 
	.data(), 
	.rden(1'b1), 
	.wren(1'b0), 
	.q(pos_data[3*DATA_WIDTH-1:2*DATA_WIDTH])
);
cell_2_3_2
#(
	.DATA_WIDTH(DATA_WIDTH), 
	.PARTICLE_NUM(PARTICLE_NUM), 
	.ADDR_WIDTH(7)
)
pos_cache_2_3_2
(
	.address(particle_id), 
	.clock(clk), 
	.data(), 
	.rden(1'b1), 
	.wren(1'b0), 
	.q(pos_data[4*DATA_WIDTH-1:3*DATA_WIDTH])
);
cell_2_3_3
#(
	.DATA_WIDTH(DATA_WIDTH), 
	.PARTICLE_NUM(PARTICLE_NUM), 
	.ADDR_WIDTH(7)
)
pos_cache_2_3_3
(
	.address(particle_id), 
	.clock(clk), 
	.data(), 
	.rden(1'b1), 
	.wren(1'b0), 
	.q(pos_data[5*DATA_WIDTH-1:4*DATA_WIDTH])
);
cell_3_1_1
#(
	.DATA_WIDTH(DATA_WIDTH), 
	.PARTICLE_NUM(PARTICLE_NUM), 
	.ADDR_WIDTH(7)
)
pos_cache_3_1_1
(
	.address(particle_id), 
	.clock(clk), 
	.data(), 
	.rden(1'b1), 
	.wren(1'b0), 
	.q(pos_data[6*DATA_WIDTH-1:5*DATA_WIDTH])
);
cell_3_1_2
#(
	.DATA_WIDTH(DATA_WIDTH), 
	.PARTICLE_NUM(PARTICLE_NUM), 
	.ADDR_WIDTH(7)
)
pos_cache_3_1_2
(
	.address(particle_id), 
	.clock(clk), 
	.data(), 
	.rden(1'b1), 
	.wren(1'b0), 
	.q(pos_data[7*DATA_WIDTH-1:6*DATA_WIDTH])
);
cell_3_1_3
#(
	.DATA_WIDTH(DATA_WIDTH), 
	.PARTICLE_NUM(PARTICLE_NUM), 
	.ADDR_WIDTH(7)
)
pos_cache_3_1_3
(
	.address(particle_id), 
	.clock(clk), 
	.data(), 
	.rden(1'b1), 
	.wren(1'b0), 
	.q(pos_data[8*DATA_WIDTH-1:7*DATA_WIDTH])
);
cell_3_2_1
#(
	.DATA_WIDTH(DATA_WIDTH), 
	.PARTICLE_NUM(PARTICLE_NUM), 
	.ADDR_WIDTH(7)
)
pos_cache_3_2_1
(
	.address(particle_id), 
	.clock(clk), 
	.data(), 
	.rden(1'b1), 
	.wren(1'b0), 
	.q(pos_data[9*DATA_WIDTH-1:8*DATA_WIDTH])
);
cell_3_2_2
#(
	.DATA_WIDTH(DATA_WIDTH), 
	.PARTICLE_NUM(PARTICLE_NUM), 
	.ADDR_WIDTH(7)
)
pos_cache_3_2_2
(
	.address(particle_id), 
	.clock(clk), 
	.data(), 
	.rden(1'b1), 
	.wren(1'b0), 
	.q(pos_data[10*DATA_WIDTH-1:9*DATA_WIDTH])
);
cell_3_2_3
#(
	.DATA_WIDTH(DATA_WIDTH), 
	.PARTICLE_NUM(PARTICLE_NUM), 
	.ADDR_WIDTH(7)
)
pos_cache_3_2_3
(
	.address(particle_id), 
	.clock(clk), 
	.data(), 
	.rden(1'b1), 
	.wren(1'b0), 
	.q(pos_data[11*DATA_WIDTH-1:10*DATA_WIDTH])
);
cell_3_3_1
#(
	.DATA_WIDTH(DATA_WIDTH), 
	.PARTICLE_NUM(PARTICLE_NUM), 
	.ADDR_WIDTH(7)
)
pos_cache_3_3_1
(
	.address(particle_id), 
	.clock(clk), 
	.data(), 
	.rden(1'b1), 
	.wren(1'b0), 
	.q(pos_data[12*DATA_WIDTH-1:11*DATA_WIDTH])
);
cell_3_3_2
#(
	.DATA_WIDTH(DATA_WIDTH), 
	.PARTICLE_NUM(PARTICLE_NUM), 
	.ADDR_WIDTH(7)
)
pos_cache_3_3_2
(
	.address(particle_id), 
	.clock(clk), 
	.data(), 
	.rden(1'b1), 
	.wren(1'b0), 
	.q(pos_data[13*DATA_WIDTH-1:12*DATA_WIDTH])
);
cell_3_3_3
#(
	.DATA_WIDTH(DATA_WIDTH), 
	.PARTICLE_NUM(PARTICLE_NUM), 
	.ADDR_WIDTH(7)
)
pos_cache_3_3_3
(
	.address(particle_id), 
	.clock(clk), 
	.data(), 
	.rden(1'b1), 
	.wren(1'b0), 
	.q(pos_data[14*DATA_WIDTH-1:13*DATA_WIDTH])
);
endmodule