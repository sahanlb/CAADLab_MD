// RAM_DualPort.v

// Generated using ACDS version 18.0 219

`timescale 1 ps / 1 ps
module RAM_DualPort (
		input  wire [12287:0] data,      //  ram_input.datain
		input  wire [4:0]     wraddress, //           .wraddress
		input  wire [9:0]     rdaddress, //           .rdaddress
		input  wire           wren,      //           .wren
		input  wire           clock,     //           .clock
		output wire [383:0]   q          // ram_output.dataout
	);

	RAM_DualPort_ram_2port_180_l4n36dy ram_2port_0 (
		.data      (data),      //   input,  width = 12288,  ram_input.datain
		.wraddress (wraddress), //   input,      width = 5,           .wraddress
		.rdaddress (rdaddress), //   input,     width = 10,           .rdaddress
		.wren      (wren),      //   input,      width = 1,           .wren
		.clock     (clock),     //   input,      width = 1,           .clock
		.q         (q)          //  output,    width = 384, ram_output.dataout
	);

endmodule
