`include "define.v"

module all_velocity_caches
#(
	parameter NUM_CELLS = 64, 
	parameter DATA_WIDTH = 32, 
	parameter CELL_ID_WIDTH = 3,
	parameter NUM_PARTICLE_PER_CELL = 128, 
	parameter PARTICLE_ID_WIDTH = 7
)
(
	input clk,
	input rst,
	input Motion_Update_enable,
	input [PARTICLE_ID_WIDTH-1:0] MU_rd_addr,
	input [3*DATA_WIDTH-1:0] MU_wr_data,
	input [3*CELL_ID_WIDTH-1:0] MU_dst_cell,
	input MU_wr_data_valid,
	input MU_rden,
	
	output [NUM_CELLS-1:0][*3*DATA_WIDTH-1:0] velocity_data_out
);

`VELOCITY_CACHE_INSTANCE(1,1,1)
`VELOCITY_CACHE_INSTANCE(1,1,2)
`VELOCITY_CACHE_INSTANCE(1,1,3)
`VELOCITY_CACHE_INSTANCE(1,1,4)
`VELOCITY_CACHE_INSTANCE(1,1,5)
`VELOCITY_CACHE_INSTANCE(1,2,1)
`VELOCITY_CACHE_INSTANCE(1,2,2)
`VELOCITY_CACHE_INSTANCE(1,2,3)
`VELOCITY_CACHE_INSTANCE(1,2,4)
`VELOCITY_CACHE_INSTANCE(1,2,5)
`VELOCITY_CACHE_INSTANCE(1,3,1)
`VELOCITY_CACHE_INSTANCE(1,3,2)
`VELOCITY_CACHE_INSTANCE(1,3,3)
`VELOCITY_CACHE_INSTANCE(1,3,4)
`VELOCITY_CACHE_INSTANCE(1,3,5)
`VELOCITY_CACHE_INSTANCE(1,4,1)
`VELOCITY_CACHE_INSTANCE(1,4,2)
`VELOCITY_CACHE_INSTANCE(1,4,3)
`VELOCITY_CACHE_INSTANCE(1,4,4)
`VELOCITY_CACHE_INSTANCE(1,4,5)
`VELOCITY_CACHE_INSTANCE(1,5,1)
`VELOCITY_CACHE_INSTANCE(1,5,2)
`VELOCITY_CACHE_INSTANCE(1,5,3)
`VELOCITY_CACHE_INSTANCE(1,5,4)
`VELOCITY_CACHE_INSTANCE(1,5,5)
`VELOCITY_CACHE_INSTANCE(2,1,1)
`VELOCITY_CACHE_INSTANCE(2,1,2)
`VELOCITY_CACHE_INSTANCE(2,1,3)
`VELOCITY_CACHE_INSTANCE(2,1,4)
`VELOCITY_CACHE_INSTANCE(2,1,5)
`VELOCITY_CACHE_INSTANCE(2,2,1)
`VELOCITY_CACHE_INSTANCE(2,2,2)
`VELOCITY_CACHE_INSTANCE(2,2,3)
`VELOCITY_CACHE_INSTANCE(2,2,4)
`VELOCITY_CACHE_INSTANCE(2,2,5)
`VELOCITY_CACHE_INSTANCE(2,3,1)
`VELOCITY_CACHE_INSTANCE(2,3,2)
`VELOCITY_CACHE_INSTANCE(2,3,3)
`VELOCITY_CACHE_INSTANCE(2,3,4)
`VELOCITY_CACHE_INSTANCE(2,3,5)
`VELOCITY_CACHE_INSTANCE(2,4,1)
`VELOCITY_CACHE_INSTANCE(2,4,2)
`VELOCITY_CACHE_INSTANCE(2,4,3)
`VELOCITY_CACHE_INSTANCE(2,4,4)
`VELOCITY_CACHE_INSTANCE(2,4,5)
`VELOCITY_CACHE_INSTANCE(2,5,1)
`VELOCITY_CACHE_INSTANCE(2,5,2)
`VELOCITY_CACHE_INSTANCE(2,5,3)
`VELOCITY_CACHE_INSTANCE(2,5,4)
`VELOCITY_CACHE_INSTANCE(2,5,5)
`VELOCITY_CACHE_INSTANCE(3,1,1)
`VELOCITY_CACHE_INSTANCE(3,1,2)
`VELOCITY_CACHE_INSTANCE(3,1,3)
`VELOCITY_CACHE_INSTANCE(3,1,4)
`VELOCITY_CACHE_INSTANCE(3,1,5)
`VELOCITY_CACHE_INSTANCE(3,2,1)
`VELOCITY_CACHE_INSTANCE(3,2,2)
`VELOCITY_CACHE_INSTANCE(3,2,3)
`VELOCITY_CACHE_INSTANCE(3,2,4)
`VELOCITY_CACHE_INSTANCE(3,2,5)
`VELOCITY_CACHE_INSTANCE(3,3,1)
`VELOCITY_CACHE_INSTANCE(3,3,2)
`VELOCITY_CACHE_INSTANCE(3,3,3)
`VELOCITY_CACHE_INSTANCE(3,3,4)
`VELOCITY_CACHE_INSTANCE(3,3,5)
`VELOCITY_CACHE_INSTANCE(3,4,1)
`VELOCITY_CACHE_INSTANCE(3,4,2)
`VELOCITY_CACHE_INSTANCE(3,4,3)
`VELOCITY_CACHE_INSTANCE(3,4,4)
`VELOCITY_CACHE_INSTANCE(3,4,5)
`VELOCITY_CACHE_INSTANCE(3,5,1)
`VELOCITY_CACHE_INSTANCE(3,5,2)
`VELOCITY_CACHE_INSTANCE(3,5,3)
`VELOCITY_CACHE_INSTANCE(3,5,4)
`VELOCITY_CACHE_INSTANCE(3,5,5)
`VELOCITY_CACHE_INSTANCE(4,1,1)
`VELOCITY_CACHE_INSTANCE(4,1,2)
`VELOCITY_CACHE_INSTANCE(4,1,3)
`VELOCITY_CACHE_INSTANCE(4,1,4)
`VELOCITY_CACHE_INSTANCE(4,1,5)
`VELOCITY_CACHE_INSTANCE(4,2,1)
`VELOCITY_CACHE_INSTANCE(4,2,2)
`VELOCITY_CACHE_INSTANCE(4,2,3)
`VELOCITY_CACHE_INSTANCE(4,2,4)
`VELOCITY_CACHE_INSTANCE(4,2,5)
`VELOCITY_CACHE_INSTANCE(4,3,1)
`VELOCITY_CACHE_INSTANCE(4,3,2)
`VELOCITY_CACHE_INSTANCE(4,3,3)
`VELOCITY_CACHE_INSTANCE(4,3,4)
`VELOCITY_CACHE_INSTANCE(4,3,5)
`VELOCITY_CACHE_INSTANCE(4,4,1)
`VELOCITY_CACHE_INSTANCE(4,4,2)
`VELOCITY_CACHE_INSTANCE(4,4,3)
`VELOCITY_CACHE_INSTANCE(4,4,4)
`VELOCITY_CACHE_INSTANCE(4,4,5)
`VELOCITY_CACHE_INSTANCE(4,5,1)
`VELOCITY_CACHE_INSTANCE(4,5,2)
`VELOCITY_CACHE_INSTANCE(4,5,3)
`VELOCITY_CACHE_INSTANCE(4,5,4)
`VELOCITY_CACHE_INSTANCE(4,5,5)
`VELOCITY_CACHE_INSTANCE(5,1,1)
`VELOCITY_CACHE_INSTANCE(5,1,2)
`VELOCITY_CACHE_INSTANCE(5,1,3)
`VELOCITY_CACHE_INSTANCE(5,1,4)
`VELOCITY_CACHE_INSTANCE(5,1,5)
`VELOCITY_CACHE_INSTANCE(5,2,1)
`VELOCITY_CACHE_INSTANCE(5,2,2)
`VELOCITY_CACHE_INSTANCE(5,2,3)
`VELOCITY_CACHE_INSTANCE(5,2,4)
`VELOCITY_CACHE_INSTANCE(5,2,5)
`VELOCITY_CACHE_INSTANCE(5,3,1)
`VELOCITY_CACHE_INSTANCE(5,3,2)
`VELOCITY_CACHE_INSTANCE(5,3,3)
`VELOCITY_CACHE_INSTANCE(5,3,4)
`VELOCITY_CACHE_INSTANCE(5,3,5)
`VELOCITY_CACHE_INSTANCE(5,4,1)
`VELOCITY_CACHE_INSTANCE(5,4,2)
`VELOCITY_CACHE_INSTANCE(5,4,3)
`VELOCITY_CACHE_INSTANCE(5,4,4)
`VELOCITY_CACHE_INSTANCE(5,4,5)
`VELOCITY_CACHE_INSTANCE(5,5,1)
`VELOCITY_CACHE_INSTANCE(5,5,2)
`VELOCITY_CACHE_INSTANCE(5,5,3)
`VELOCITY_CACHE_INSTANCE(5,5,4)
`VELOCITY_CACHE_INSTANCE(5,5,5)
	
endmodule
