module FIX_ADD (
		input  wire [31:0] a0,     //     a0.a0
		input  wire [31:0] a1,     //     a1.a1
		input  wire        clk,    //    clk.clk
		input  wire [0:0]  en,     //     en.en
		output wire [31:0] result, // result.result
		input  wire        rst     //    rst.reset
	);
endmodule

