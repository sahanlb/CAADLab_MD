// Int_Mul_Add.v

// Generated using ACDS version 18.0 219

`timescale 1 ps / 1 ps
module Int_Mul_Add (
		input  wire [3:0] dataa_0, // dataa_0.dataa_0
		input  wire [3:0] datab_0, // datab_0.datab_0
		output wire [3:0] result   //  result.result
	);

	Int_Mul_Add_altera_mult_add_180_7hdzzqq mult_add_0 (
		.result  (result),  //  output,  width = 4,  result.result
		.dataa_0 (dataa_0), //   input,  width = 4, dataa_0.dataa_0
		.datab_0 (datab_0)  //   input,  width = 4, datab_0.datab_0
	);

endmodule
