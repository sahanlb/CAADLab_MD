module FP_Sqrt (
		input  wire [31:0] a,      //      a.a
		input  wire        areset, // areset.reset
		input  wire        clk,    //    clk.clk
		output wire [31:0] q       //      q.q
	);
endmodule

