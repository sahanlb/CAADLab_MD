module FIX_MUL (
		input  wire [31:0] a,      //      a.a
		input  wire [31:0] b,      //      b.b
		input  wire        clk,    //    clk.clk
		input  wire [0:0]  en,     //     en.en
		output wire [63:0] result, // result.result
		input  wire        rst     //    rst.reset
	);
endmodule

