// FIFO2.v

// Generated using ACDS version 18.0 219

`timescale 1 ps / 1 ps
module filter_buffer_MLAB 
	#(
		parameter FILTER_BUFFER_DATA_WIDTH = 224
	)
	(
		input  wire [FILTER_BUFFER_DATA_WIDTH-1:0] w_data,  //  fifo2_input.w_data
		input  wire         w_req,   //             .w_req
		input  wire         r_req,   //             .r_req
		input  wire         clk,     //             .clk
		input  wire         sclr,    //             .sclr
		output wire [FILTER_BUFFER_DATA_WIDTH-1:0] r_data,  // fifo2_output.r_data
		output wire [4:0]   w_usedw, //             .w_usedw
		output wire [4:0]   r_usedw, //             .r_usedw
		output wire         w_full,  //             .w_full
		output wire         w_ready, //             .w_ready
		output wire         r_empty, //             .r_empty
		output wire         r_valid  //             .r_valid
	);

	FIFO2_fifo2_180_bd2zssi #(
		.SCFIFO_MODE         (1),
		.DATAWIDTH           (FILTER_BUFFER_DATA_WIDTH),
		.RAM_BLK_TYPE        ("MLAB"),
		.USE_ACLR_PORT       (0),
		.RAM_WRPTR_DUPLICATE (0),
		.RAM_RDPTR_DUPLICATE (0)
	) fifo2_0 (
		.w_data  (w_data),  //   input,  width = 200,  fifo2_input.w_data
		.w_req   (w_req),   //   input,    width = 1,             .w_req
		.r_req   (r_req),   //   input,    width = 1,             .r_req
		.clk     (clk),     //   input,    width = 1,             .clk
		.sclr    (sclr),    //   input,    width = 1,             .sclr
		.r_data  (r_data),  //  output,  width = 200, fifo2_output.r_data
		.w_usedw (w_usedw), //  output,    width = 5,             .w_usedw
		.r_usedw (r_usedw), //  output,    width = 5,             .r_usedw
		.w_full  (w_full),  //  output,    width = 1,             .w_full
		.w_ready (w_ready), //  output,    width = 1,             .w_ready
		.r_empty (r_empty), //  output,    width = 1,             .r_empty
		.r_valid (r_valid), //  output,    width = 1,             .r_valid
		.aclr    (1'b0),    // (terminated),                            
		.w_clk   (1'b0),    // (terminated),                            
		.r_clk   (1'b0),    // (terminated),                            
		.w_sclr  (1'b0),    // (terminated),                            
		.r_sclr  (1'b0),    // (terminated),                            
		.w_aclr  (1'b0),    // (terminated),                            
		.r_aclr  (1'b0)     // (terminated),                            
	);

endmodule
