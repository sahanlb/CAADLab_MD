// FP_GreaterThan_or_Equal.v

// Generated using ACDS version 18.0 219

`timescale 1 ps / 1 ps
module FP_GreaterThan_or_Equal (
		input  wire [31:0] a,      //      a.a
		input  wire        areset, // areset.reset
		input  wire [31:0] b,      //      b.b
		input  wire        clk,    //    clk.clk
		output wire [0:0]  q       //      q.q
	);

	FP_GreaterThan_or_Equal_altera_fp_functions_180_nqpmigq fp_functions_0 (
		.clk    (clk),    //   input,   width = 1,    clk.clk
		.areset (areset), //   input,   width = 1, areset.reset
		.a      (a),      //   input,  width = 32,      a.a
		.b      (b),      //   input,  width = 32,      b.b
		.q      (q)       //  output,   width = 1,      q.q
	);

endmodule
