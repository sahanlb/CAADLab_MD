module force_to_valid_force_mapping
#(
	parameter DATA_WIDTH = 32, 
	parameter NUM_CELLS = 64, 
	parameter NUM_NEIGHBOR_CELLS = 13, 
	parameter NUM_FILTER = 7, 
	parameter PARTICLE_ID_WIDTH = 7, 
	parameter FORCE_BUFFER_WIDTH = 3*DATA_WIDTH+PARTICLE_ID_WIDTH+1, 
	parameter FORCE_DATA_WIDTH = FORCE_BUFFER_WIDTH-1
)
(
	input [NUM_CELLS*(NUM_NEIGHBOR_CELLS+1)-1:0] arbitration_result, 
	input [NUM_CELLS*NUM_FILTER*FORCE_DATA_WIDTH-1:0] force_and_addr, 
	
	output reg [NUM_CELLS*FORCE_DATA_WIDTH-1:0] force_to_caches
);

always@(*)
	begin
	case(arbitration_result[1*(NUM_NEIGHBOR_CELLS+1)-1:0*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[1*FORCE_DATA_WIDTH-1:0*FORCE_DATA_WIDTH] = force_and_addr[0*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:0*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[1*FORCE_DATA_WIDTH-1:0*FORCE_DATA_WIDTH] = force_and_addr[3*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:3*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[1*FORCE_DATA_WIDTH-1:0*FORCE_DATA_WIDTH] = force_and_addr[4*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:4*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[1*FORCE_DATA_WIDTH-1:0*FORCE_DATA_WIDTH] = force_and_addr[5*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:5*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[1*FORCE_DATA_WIDTH-1:0*FORCE_DATA_WIDTH] = force_and_addr[13*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:13*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[1*FORCE_DATA_WIDTH-1:0*FORCE_DATA_WIDTH] = force_and_addr[17*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:17*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[1*FORCE_DATA_WIDTH-1:0*FORCE_DATA_WIDTH] = force_and_addr[19*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:19*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[1*FORCE_DATA_WIDTH-1:0*FORCE_DATA_WIDTH] = force_and_addr[21*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:21*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[1*FORCE_DATA_WIDTH-1:0*FORCE_DATA_WIDTH] = force_and_addr[28*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:28*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[1*FORCE_DATA_WIDTH-1:0*FORCE_DATA_WIDTH] = force_and_addr[29*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:29*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[1*FORCE_DATA_WIDTH-1:0*FORCE_DATA_WIDTH] = force_and_addr[48*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:48*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[1*FORCE_DATA_WIDTH-1:0*FORCE_DATA_WIDTH] = force_and_addr[53*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:53*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[1*FORCE_DATA_WIDTH-1:0*FORCE_DATA_WIDTH] = force_and_addr[60*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:60*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[1*FORCE_DATA_WIDTH-1:0*FORCE_DATA_WIDTH] = force_and_addr[61*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:61*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[1*FORCE_DATA_WIDTH-1:0*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[2*(NUM_NEIGHBOR_CELLS+1)-1:1*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[2*FORCE_DATA_WIDTH-1:1*FORCE_DATA_WIDTH] = force_and_addr[0*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:0*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[2*FORCE_DATA_WIDTH-1:1*FORCE_DATA_WIDTH] = force_and_addr[1*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:1*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[2*FORCE_DATA_WIDTH-1:1*FORCE_DATA_WIDTH] = force_and_addr[5*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:5*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[2*FORCE_DATA_WIDTH-1:1*FORCE_DATA_WIDTH] = force_and_addr[6*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:6*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[2*FORCE_DATA_WIDTH-1:1*FORCE_DATA_WIDTH] = force_and_addr[14*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:14*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[2*FORCE_DATA_WIDTH-1:1*FORCE_DATA_WIDTH] = force_and_addr[16*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:16*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[2*FORCE_DATA_WIDTH-1:1*FORCE_DATA_WIDTH] = force_and_addr[18*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:18*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[2*FORCE_DATA_WIDTH-1:1*FORCE_DATA_WIDTH] = force_and_addr[22*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:22*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[2*FORCE_DATA_WIDTH-1:1*FORCE_DATA_WIDTH] = force_and_addr[29*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:29*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[2*FORCE_DATA_WIDTH-1:1*FORCE_DATA_WIDTH] = force_and_addr[30*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:30*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[2*FORCE_DATA_WIDTH-1:1*FORCE_DATA_WIDTH] = force_and_addr[49*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:49*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[2*FORCE_DATA_WIDTH-1:1*FORCE_DATA_WIDTH] = force_and_addr[54*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:54*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[2*FORCE_DATA_WIDTH-1:1*FORCE_DATA_WIDTH] = force_and_addr[61*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:61*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[2*FORCE_DATA_WIDTH-1:1*FORCE_DATA_WIDTH] = force_and_addr[62*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:62*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[2*FORCE_DATA_WIDTH-1:1*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[3*(NUM_NEIGHBOR_CELLS+1)-1:2*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[3*FORCE_DATA_WIDTH-1:2*FORCE_DATA_WIDTH] = force_and_addr[1*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:1*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[3*FORCE_DATA_WIDTH-1:2*FORCE_DATA_WIDTH] = force_and_addr[2*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:2*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[3*FORCE_DATA_WIDTH-1:2*FORCE_DATA_WIDTH] = force_and_addr[6*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:6*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[3*FORCE_DATA_WIDTH-1:2*FORCE_DATA_WIDTH] = force_and_addr[7*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:7*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[3*FORCE_DATA_WIDTH-1:2*FORCE_DATA_WIDTH] = force_and_addr[15*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:15*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[3*FORCE_DATA_WIDTH-1:2*FORCE_DATA_WIDTH] = force_and_addr[17*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:17*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[3*FORCE_DATA_WIDTH-1:2*FORCE_DATA_WIDTH] = force_and_addr[19*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:19*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[3*FORCE_DATA_WIDTH-1:2*FORCE_DATA_WIDTH] = force_and_addr[23*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:23*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[3*FORCE_DATA_WIDTH-1:2*FORCE_DATA_WIDTH] = force_and_addr[30*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:30*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[3*FORCE_DATA_WIDTH-1:2*FORCE_DATA_WIDTH] = force_and_addr[31*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:31*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[3*FORCE_DATA_WIDTH-1:2*FORCE_DATA_WIDTH] = force_and_addr[50*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:50*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[3*FORCE_DATA_WIDTH-1:2*FORCE_DATA_WIDTH] = force_and_addr[55*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:55*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[3*FORCE_DATA_WIDTH-1:2*FORCE_DATA_WIDTH] = force_and_addr[62*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:62*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[3*FORCE_DATA_WIDTH-1:2*FORCE_DATA_WIDTH] = force_and_addr[63*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:63*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[3*FORCE_DATA_WIDTH-1:2*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[4*(NUM_NEIGHBOR_CELLS+1)-1:3*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[4*FORCE_DATA_WIDTH-1:3*FORCE_DATA_WIDTH] = force_and_addr[2*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:2*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[4*FORCE_DATA_WIDTH-1:3*FORCE_DATA_WIDTH] = force_and_addr[3*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:3*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[4*FORCE_DATA_WIDTH-1:3*FORCE_DATA_WIDTH] = force_and_addr[4*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:4*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[4*FORCE_DATA_WIDTH-1:3*FORCE_DATA_WIDTH] = force_and_addr[7*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:7*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[4*FORCE_DATA_WIDTH-1:3*FORCE_DATA_WIDTH] = force_and_addr[12*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:12*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[4*FORCE_DATA_WIDTH-1:3*FORCE_DATA_WIDTH] = force_and_addr[16*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:16*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[4*FORCE_DATA_WIDTH-1:3*FORCE_DATA_WIDTH] = force_and_addr[18*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:18*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[4*FORCE_DATA_WIDTH-1:3*FORCE_DATA_WIDTH] = force_and_addr[20*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:20*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[4*FORCE_DATA_WIDTH-1:3*FORCE_DATA_WIDTH] = force_and_addr[28*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:28*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[4*FORCE_DATA_WIDTH-1:3*FORCE_DATA_WIDTH] = force_and_addr[31*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:31*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[4*FORCE_DATA_WIDTH-1:3*FORCE_DATA_WIDTH] = force_and_addr[51*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:51*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[4*FORCE_DATA_WIDTH-1:3*FORCE_DATA_WIDTH] = force_and_addr[52*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:52*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[4*FORCE_DATA_WIDTH-1:3*FORCE_DATA_WIDTH] = force_and_addr[60*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:60*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[4*FORCE_DATA_WIDTH-1:3*FORCE_DATA_WIDTH] = force_and_addr[63*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:63*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[4*FORCE_DATA_WIDTH-1:3*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[5*(NUM_NEIGHBOR_CELLS+1)-1:4*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[5*FORCE_DATA_WIDTH-1:4*FORCE_DATA_WIDTH] = force_and_addr[1*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:1*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[5*FORCE_DATA_WIDTH-1:4*FORCE_DATA_WIDTH] = force_and_addr[4*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:4*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[5*FORCE_DATA_WIDTH-1:4*FORCE_DATA_WIDTH] = force_and_addr[7*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:7*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[5*FORCE_DATA_WIDTH-1:4*FORCE_DATA_WIDTH] = force_and_addr[8*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:8*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[5*FORCE_DATA_WIDTH-1:4*FORCE_DATA_WIDTH] = force_and_addr[9*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:9*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[5*FORCE_DATA_WIDTH-1:4*FORCE_DATA_WIDTH] = force_and_addr[16*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:16*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[5*FORCE_DATA_WIDTH-1:4*FORCE_DATA_WIDTH] = force_and_addr[17*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:17*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[5*FORCE_DATA_WIDTH-1:4*FORCE_DATA_WIDTH] = force_and_addr[21*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:21*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[5*FORCE_DATA_WIDTH-1:4*FORCE_DATA_WIDTH] = force_and_addr[23*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:23*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[5*FORCE_DATA_WIDTH-1:4*FORCE_DATA_WIDTH] = force_and_addr[25*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:25*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[5*FORCE_DATA_WIDTH-1:4*FORCE_DATA_WIDTH] = force_and_addr[48*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:48*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[5*FORCE_DATA_WIDTH-1:4*FORCE_DATA_WIDTH] = force_and_addr[49*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:49*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[5*FORCE_DATA_WIDTH-1:4*FORCE_DATA_WIDTH] = force_and_addr[52*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:52*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[5*FORCE_DATA_WIDTH-1:4*FORCE_DATA_WIDTH] = force_and_addr[57*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:57*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[5*FORCE_DATA_WIDTH-1:4*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[6*(NUM_NEIGHBOR_CELLS+1)-1:5*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[6*FORCE_DATA_WIDTH-1:5*FORCE_DATA_WIDTH] = force_and_addr[2*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:2*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[6*FORCE_DATA_WIDTH-1:5*FORCE_DATA_WIDTH] = force_and_addr[4*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:4*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[6*FORCE_DATA_WIDTH-1:5*FORCE_DATA_WIDTH] = force_and_addr[5*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:5*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[6*FORCE_DATA_WIDTH-1:5*FORCE_DATA_WIDTH] = force_and_addr[9*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:9*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[6*FORCE_DATA_WIDTH-1:5*FORCE_DATA_WIDTH] = force_and_addr[10*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:10*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[6*FORCE_DATA_WIDTH-1:5*FORCE_DATA_WIDTH] = force_and_addr[17*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:17*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[6*FORCE_DATA_WIDTH-1:5*FORCE_DATA_WIDTH] = force_and_addr[18*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:18*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[6*FORCE_DATA_WIDTH-1:5*FORCE_DATA_WIDTH] = force_and_addr[20*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:20*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[6*FORCE_DATA_WIDTH-1:5*FORCE_DATA_WIDTH] = force_and_addr[22*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:22*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[6*FORCE_DATA_WIDTH-1:5*FORCE_DATA_WIDTH] = force_and_addr[26*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:26*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[6*FORCE_DATA_WIDTH-1:5*FORCE_DATA_WIDTH] = force_and_addr[49*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:49*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[6*FORCE_DATA_WIDTH-1:5*FORCE_DATA_WIDTH] = force_and_addr[50*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:50*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[6*FORCE_DATA_WIDTH-1:5*FORCE_DATA_WIDTH] = force_and_addr[53*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:53*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[6*FORCE_DATA_WIDTH-1:5*FORCE_DATA_WIDTH] = force_and_addr[58*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:58*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[6*FORCE_DATA_WIDTH-1:5*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[7*(NUM_NEIGHBOR_CELLS+1)-1:6*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[7*FORCE_DATA_WIDTH-1:6*FORCE_DATA_WIDTH] = force_and_addr[3*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:3*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[7*FORCE_DATA_WIDTH-1:6*FORCE_DATA_WIDTH] = force_and_addr[5*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:5*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[7*FORCE_DATA_WIDTH-1:6*FORCE_DATA_WIDTH] = force_and_addr[6*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:6*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[7*FORCE_DATA_WIDTH-1:6*FORCE_DATA_WIDTH] = force_and_addr[10*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:10*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[7*FORCE_DATA_WIDTH-1:6*FORCE_DATA_WIDTH] = force_and_addr[11*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:11*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[7*FORCE_DATA_WIDTH-1:6*FORCE_DATA_WIDTH] = force_and_addr[18*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:18*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[7*FORCE_DATA_WIDTH-1:6*FORCE_DATA_WIDTH] = force_and_addr[19*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:19*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[7*FORCE_DATA_WIDTH-1:6*FORCE_DATA_WIDTH] = force_and_addr[21*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:21*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[7*FORCE_DATA_WIDTH-1:6*FORCE_DATA_WIDTH] = force_and_addr[23*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:23*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[7*FORCE_DATA_WIDTH-1:6*FORCE_DATA_WIDTH] = force_and_addr[27*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:27*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[7*FORCE_DATA_WIDTH-1:6*FORCE_DATA_WIDTH] = force_and_addr[50*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:50*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[7*FORCE_DATA_WIDTH-1:6*FORCE_DATA_WIDTH] = force_and_addr[51*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:51*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[7*FORCE_DATA_WIDTH-1:6*FORCE_DATA_WIDTH] = force_and_addr[54*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:54*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[7*FORCE_DATA_WIDTH-1:6*FORCE_DATA_WIDTH] = force_and_addr[59*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:59*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[7*FORCE_DATA_WIDTH-1:6*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[8*(NUM_NEIGHBOR_CELLS+1)-1:7*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[8*FORCE_DATA_WIDTH-1:7*FORCE_DATA_WIDTH] = force_and_addr[0*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:0*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[8*FORCE_DATA_WIDTH-1:7*FORCE_DATA_WIDTH] = force_and_addr[6*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:6*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[8*FORCE_DATA_WIDTH-1:7*FORCE_DATA_WIDTH] = force_and_addr[7*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:7*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[8*FORCE_DATA_WIDTH-1:7*FORCE_DATA_WIDTH] = force_and_addr[8*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:8*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[8*FORCE_DATA_WIDTH-1:7*FORCE_DATA_WIDTH] = force_and_addr[11*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:11*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[8*FORCE_DATA_WIDTH-1:7*FORCE_DATA_WIDTH] = force_and_addr[16*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:16*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[8*FORCE_DATA_WIDTH-1:7*FORCE_DATA_WIDTH] = force_and_addr[19*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:19*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[8*FORCE_DATA_WIDTH-1:7*FORCE_DATA_WIDTH] = force_and_addr[20*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:20*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[8*FORCE_DATA_WIDTH-1:7*FORCE_DATA_WIDTH] = force_and_addr[22*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:22*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[8*FORCE_DATA_WIDTH-1:7*FORCE_DATA_WIDTH] = force_and_addr[24*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:24*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[8*FORCE_DATA_WIDTH-1:7*FORCE_DATA_WIDTH] = force_and_addr[48*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:48*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[8*FORCE_DATA_WIDTH-1:7*FORCE_DATA_WIDTH] = force_and_addr[51*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:51*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[8*FORCE_DATA_WIDTH-1:7*FORCE_DATA_WIDTH] = force_and_addr[55*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:55*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[8*FORCE_DATA_WIDTH-1:7*FORCE_DATA_WIDTH] = force_and_addr[56*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:56*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[8*FORCE_DATA_WIDTH-1:7*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[9*(NUM_NEIGHBOR_CELLS+1)-1:8*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[9*FORCE_DATA_WIDTH-1:8*FORCE_DATA_WIDTH] = force_and_addr[5*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:5*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[9*FORCE_DATA_WIDTH-1:8*FORCE_DATA_WIDTH] = force_and_addr[8*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:8*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[9*FORCE_DATA_WIDTH-1:8*FORCE_DATA_WIDTH] = force_and_addr[11*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:11*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[9*FORCE_DATA_WIDTH-1:8*FORCE_DATA_WIDTH] = force_and_addr[12*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:12*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[9*FORCE_DATA_WIDTH-1:8*FORCE_DATA_WIDTH] = force_and_addr[13*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:13*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[9*FORCE_DATA_WIDTH-1:8*FORCE_DATA_WIDTH] = force_and_addr[20*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:20*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[9*FORCE_DATA_WIDTH-1:8*FORCE_DATA_WIDTH] = force_and_addr[21*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:21*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[9*FORCE_DATA_WIDTH-1:8*FORCE_DATA_WIDTH] = force_and_addr[25*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:25*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[9*FORCE_DATA_WIDTH-1:8*FORCE_DATA_WIDTH] = force_and_addr[27*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:27*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[9*FORCE_DATA_WIDTH-1:8*FORCE_DATA_WIDTH] = force_and_addr[29*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:29*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[9*FORCE_DATA_WIDTH-1:8*FORCE_DATA_WIDTH] = force_and_addr[52*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:52*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[9*FORCE_DATA_WIDTH-1:8*FORCE_DATA_WIDTH] = force_and_addr[53*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:53*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[9*FORCE_DATA_WIDTH-1:8*FORCE_DATA_WIDTH] = force_and_addr[56*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:56*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[9*FORCE_DATA_WIDTH-1:8*FORCE_DATA_WIDTH] = force_and_addr[61*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:61*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[9*FORCE_DATA_WIDTH-1:8*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[10*(NUM_NEIGHBOR_CELLS+1)-1:9*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[10*FORCE_DATA_WIDTH-1:9*FORCE_DATA_WIDTH] = force_and_addr[6*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:6*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[10*FORCE_DATA_WIDTH-1:9*FORCE_DATA_WIDTH] = force_and_addr[8*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:8*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[10*FORCE_DATA_WIDTH-1:9*FORCE_DATA_WIDTH] = force_and_addr[9*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:9*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[10*FORCE_DATA_WIDTH-1:9*FORCE_DATA_WIDTH] = force_and_addr[13*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:13*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[10*FORCE_DATA_WIDTH-1:9*FORCE_DATA_WIDTH] = force_and_addr[14*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:14*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[10*FORCE_DATA_WIDTH-1:9*FORCE_DATA_WIDTH] = force_and_addr[21*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:21*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[10*FORCE_DATA_WIDTH-1:9*FORCE_DATA_WIDTH] = force_and_addr[22*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:22*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[10*FORCE_DATA_WIDTH-1:9*FORCE_DATA_WIDTH] = force_and_addr[24*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:24*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[10*FORCE_DATA_WIDTH-1:9*FORCE_DATA_WIDTH] = force_and_addr[26*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:26*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[10*FORCE_DATA_WIDTH-1:9*FORCE_DATA_WIDTH] = force_and_addr[30*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:30*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[10*FORCE_DATA_WIDTH-1:9*FORCE_DATA_WIDTH] = force_and_addr[53*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:53*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[10*FORCE_DATA_WIDTH-1:9*FORCE_DATA_WIDTH] = force_and_addr[54*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:54*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[10*FORCE_DATA_WIDTH-1:9*FORCE_DATA_WIDTH] = force_and_addr[57*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:57*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[10*FORCE_DATA_WIDTH-1:9*FORCE_DATA_WIDTH] = force_and_addr[62*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:62*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[10*FORCE_DATA_WIDTH-1:9*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[11*(NUM_NEIGHBOR_CELLS+1)-1:10*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[11*FORCE_DATA_WIDTH-1:10*FORCE_DATA_WIDTH] = force_and_addr[7*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:7*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[11*FORCE_DATA_WIDTH-1:10*FORCE_DATA_WIDTH] = force_and_addr[9*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:9*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[11*FORCE_DATA_WIDTH-1:10*FORCE_DATA_WIDTH] = force_and_addr[10*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:10*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[11*FORCE_DATA_WIDTH-1:10*FORCE_DATA_WIDTH] = force_and_addr[14*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:14*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[11*FORCE_DATA_WIDTH-1:10*FORCE_DATA_WIDTH] = force_and_addr[15*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:15*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[11*FORCE_DATA_WIDTH-1:10*FORCE_DATA_WIDTH] = force_and_addr[22*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:22*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[11*FORCE_DATA_WIDTH-1:10*FORCE_DATA_WIDTH] = force_and_addr[23*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:23*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[11*FORCE_DATA_WIDTH-1:10*FORCE_DATA_WIDTH] = force_and_addr[25*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:25*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[11*FORCE_DATA_WIDTH-1:10*FORCE_DATA_WIDTH] = force_and_addr[27*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:27*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[11*FORCE_DATA_WIDTH-1:10*FORCE_DATA_WIDTH] = force_and_addr[31*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:31*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[11*FORCE_DATA_WIDTH-1:10*FORCE_DATA_WIDTH] = force_and_addr[54*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:54*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[11*FORCE_DATA_WIDTH-1:10*FORCE_DATA_WIDTH] = force_and_addr[55*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:55*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[11*FORCE_DATA_WIDTH-1:10*FORCE_DATA_WIDTH] = force_and_addr[58*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:58*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[11*FORCE_DATA_WIDTH-1:10*FORCE_DATA_WIDTH] = force_and_addr[63*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:63*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[11*FORCE_DATA_WIDTH-1:10*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[12*(NUM_NEIGHBOR_CELLS+1)-1:11*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[12*FORCE_DATA_WIDTH-1:11*FORCE_DATA_WIDTH] = force_and_addr[4*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:4*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[12*FORCE_DATA_WIDTH-1:11*FORCE_DATA_WIDTH] = force_and_addr[10*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:10*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[12*FORCE_DATA_WIDTH-1:11*FORCE_DATA_WIDTH] = force_and_addr[11*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:11*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[12*FORCE_DATA_WIDTH-1:11*FORCE_DATA_WIDTH] = force_and_addr[12*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:12*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[12*FORCE_DATA_WIDTH-1:11*FORCE_DATA_WIDTH] = force_and_addr[15*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:15*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[12*FORCE_DATA_WIDTH-1:11*FORCE_DATA_WIDTH] = force_and_addr[20*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:20*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[12*FORCE_DATA_WIDTH-1:11*FORCE_DATA_WIDTH] = force_and_addr[23*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:23*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[12*FORCE_DATA_WIDTH-1:11*FORCE_DATA_WIDTH] = force_and_addr[24*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:24*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[12*FORCE_DATA_WIDTH-1:11*FORCE_DATA_WIDTH] = force_and_addr[26*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:26*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[12*FORCE_DATA_WIDTH-1:11*FORCE_DATA_WIDTH] = force_and_addr[28*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:28*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[12*FORCE_DATA_WIDTH-1:11*FORCE_DATA_WIDTH] = force_and_addr[52*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:52*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[12*FORCE_DATA_WIDTH-1:11*FORCE_DATA_WIDTH] = force_and_addr[55*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:55*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[12*FORCE_DATA_WIDTH-1:11*FORCE_DATA_WIDTH] = force_and_addr[59*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:59*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[12*FORCE_DATA_WIDTH-1:11*FORCE_DATA_WIDTH] = force_and_addr[60*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:60*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[12*FORCE_DATA_WIDTH-1:11*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[13*(NUM_NEIGHBOR_CELLS+1)-1:12*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[13*FORCE_DATA_WIDTH-1:12*FORCE_DATA_WIDTH] = force_and_addr[0*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:0*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[13*FORCE_DATA_WIDTH-1:12*FORCE_DATA_WIDTH] = force_and_addr[1*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:1*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[13*FORCE_DATA_WIDTH-1:12*FORCE_DATA_WIDTH] = force_and_addr[9*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:9*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[13*FORCE_DATA_WIDTH-1:12*FORCE_DATA_WIDTH] = force_and_addr[12*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:12*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[13*FORCE_DATA_WIDTH-1:12*FORCE_DATA_WIDTH] = force_and_addr[15*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:15*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[13*FORCE_DATA_WIDTH-1:12*FORCE_DATA_WIDTH] = force_and_addr[17*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:17*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[13*FORCE_DATA_WIDTH-1:12*FORCE_DATA_WIDTH] = force_and_addr[24*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:24*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[13*FORCE_DATA_WIDTH-1:12*FORCE_DATA_WIDTH] = force_and_addr[25*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:25*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[13*FORCE_DATA_WIDTH-1:12*FORCE_DATA_WIDTH] = force_and_addr[29*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:29*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[13*FORCE_DATA_WIDTH-1:12*FORCE_DATA_WIDTH] = force_and_addr[31*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:31*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[13*FORCE_DATA_WIDTH-1:12*FORCE_DATA_WIDTH] = force_and_addr[49*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:49*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[13*FORCE_DATA_WIDTH-1:12*FORCE_DATA_WIDTH] = force_and_addr[56*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:56*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[13*FORCE_DATA_WIDTH-1:12*FORCE_DATA_WIDTH] = force_and_addr[57*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:57*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[13*FORCE_DATA_WIDTH-1:12*FORCE_DATA_WIDTH] = force_and_addr[60*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:60*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[13*FORCE_DATA_WIDTH-1:12*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[14*(NUM_NEIGHBOR_CELLS+1)-1:13*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[14*FORCE_DATA_WIDTH-1:13*FORCE_DATA_WIDTH] = force_and_addr[1*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:1*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[14*FORCE_DATA_WIDTH-1:13*FORCE_DATA_WIDTH] = force_and_addr[2*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:2*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[14*FORCE_DATA_WIDTH-1:13*FORCE_DATA_WIDTH] = force_and_addr[10*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:10*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[14*FORCE_DATA_WIDTH-1:13*FORCE_DATA_WIDTH] = force_and_addr[12*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:12*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[14*FORCE_DATA_WIDTH-1:13*FORCE_DATA_WIDTH] = force_and_addr[13*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:13*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[14*FORCE_DATA_WIDTH-1:13*FORCE_DATA_WIDTH] = force_and_addr[18*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:18*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[14*FORCE_DATA_WIDTH-1:13*FORCE_DATA_WIDTH] = force_and_addr[25*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:25*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[14*FORCE_DATA_WIDTH-1:13*FORCE_DATA_WIDTH] = force_and_addr[26*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:26*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[14*FORCE_DATA_WIDTH-1:13*FORCE_DATA_WIDTH] = force_and_addr[28*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:28*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[14*FORCE_DATA_WIDTH-1:13*FORCE_DATA_WIDTH] = force_and_addr[30*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:30*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[14*FORCE_DATA_WIDTH-1:13*FORCE_DATA_WIDTH] = force_and_addr[50*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:50*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[14*FORCE_DATA_WIDTH-1:13*FORCE_DATA_WIDTH] = force_and_addr[57*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:57*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[14*FORCE_DATA_WIDTH-1:13*FORCE_DATA_WIDTH] = force_and_addr[58*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:58*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[14*FORCE_DATA_WIDTH-1:13*FORCE_DATA_WIDTH] = force_and_addr[61*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:61*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[14*FORCE_DATA_WIDTH-1:13*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[15*(NUM_NEIGHBOR_CELLS+1)-1:14*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[15*FORCE_DATA_WIDTH-1:14*FORCE_DATA_WIDTH] = force_and_addr[2*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:2*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[15*FORCE_DATA_WIDTH-1:14*FORCE_DATA_WIDTH] = force_and_addr[3*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:3*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[15*FORCE_DATA_WIDTH-1:14*FORCE_DATA_WIDTH] = force_and_addr[11*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:11*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[15*FORCE_DATA_WIDTH-1:14*FORCE_DATA_WIDTH] = force_and_addr[13*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:13*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[15*FORCE_DATA_WIDTH-1:14*FORCE_DATA_WIDTH] = force_and_addr[14*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:14*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[15*FORCE_DATA_WIDTH-1:14*FORCE_DATA_WIDTH] = force_and_addr[19*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:19*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[15*FORCE_DATA_WIDTH-1:14*FORCE_DATA_WIDTH] = force_and_addr[26*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:26*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[15*FORCE_DATA_WIDTH-1:14*FORCE_DATA_WIDTH] = force_and_addr[27*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:27*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[15*FORCE_DATA_WIDTH-1:14*FORCE_DATA_WIDTH] = force_and_addr[29*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:29*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[15*FORCE_DATA_WIDTH-1:14*FORCE_DATA_WIDTH] = force_and_addr[31*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:31*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[15*FORCE_DATA_WIDTH-1:14*FORCE_DATA_WIDTH] = force_and_addr[51*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:51*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[15*FORCE_DATA_WIDTH-1:14*FORCE_DATA_WIDTH] = force_and_addr[58*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:58*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[15*FORCE_DATA_WIDTH-1:14*FORCE_DATA_WIDTH] = force_and_addr[59*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:59*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[15*FORCE_DATA_WIDTH-1:14*FORCE_DATA_WIDTH] = force_and_addr[62*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:62*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[15*FORCE_DATA_WIDTH-1:14*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[16*(NUM_NEIGHBOR_CELLS+1)-1:15*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[16*FORCE_DATA_WIDTH-1:15*FORCE_DATA_WIDTH] = force_and_addr[0*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:0*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[16*FORCE_DATA_WIDTH-1:15*FORCE_DATA_WIDTH] = force_and_addr[3*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:3*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[16*FORCE_DATA_WIDTH-1:15*FORCE_DATA_WIDTH] = force_and_addr[8*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:8*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[16*FORCE_DATA_WIDTH-1:15*FORCE_DATA_WIDTH] = force_and_addr[14*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:14*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[16*FORCE_DATA_WIDTH-1:15*FORCE_DATA_WIDTH] = force_and_addr[15*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:15*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[16*FORCE_DATA_WIDTH-1:15*FORCE_DATA_WIDTH] = force_and_addr[16*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:16*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[16*FORCE_DATA_WIDTH-1:15*FORCE_DATA_WIDTH] = force_and_addr[24*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:24*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[16*FORCE_DATA_WIDTH-1:15*FORCE_DATA_WIDTH] = force_and_addr[27*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:27*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[16*FORCE_DATA_WIDTH-1:15*FORCE_DATA_WIDTH] = force_and_addr[28*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:28*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[16*FORCE_DATA_WIDTH-1:15*FORCE_DATA_WIDTH] = force_and_addr[30*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:30*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[16*FORCE_DATA_WIDTH-1:15*FORCE_DATA_WIDTH] = force_and_addr[48*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:48*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[16*FORCE_DATA_WIDTH-1:15*FORCE_DATA_WIDTH] = force_and_addr[56*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:56*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[16*FORCE_DATA_WIDTH-1:15*FORCE_DATA_WIDTH] = force_and_addr[59*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:59*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[16*FORCE_DATA_WIDTH-1:15*FORCE_DATA_WIDTH] = force_and_addr[63*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:63*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[16*FORCE_DATA_WIDTH-1:15*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[17*(NUM_NEIGHBOR_CELLS+1)-1:16*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[17*FORCE_DATA_WIDTH-1:16*FORCE_DATA_WIDTH] = force_and_addr[0*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:0*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[17*FORCE_DATA_WIDTH-1:16*FORCE_DATA_WIDTH] = force_and_addr[5*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:5*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[17*FORCE_DATA_WIDTH-1:16*FORCE_DATA_WIDTH] = force_and_addr[12*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:12*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[17*FORCE_DATA_WIDTH-1:16*FORCE_DATA_WIDTH] = force_and_addr[13*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:13*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[17*FORCE_DATA_WIDTH-1:16*FORCE_DATA_WIDTH] = force_and_addr[16*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:16*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[17*FORCE_DATA_WIDTH-1:16*FORCE_DATA_WIDTH] = force_and_addr[19*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:19*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[17*FORCE_DATA_WIDTH-1:16*FORCE_DATA_WIDTH] = force_and_addr[20*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:20*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[17*FORCE_DATA_WIDTH-1:16*FORCE_DATA_WIDTH] = force_and_addr[21*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:21*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[17*FORCE_DATA_WIDTH-1:16*FORCE_DATA_WIDTH] = force_and_addr[29*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:29*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[17*FORCE_DATA_WIDTH-1:16*FORCE_DATA_WIDTH] = force_and_addr[33*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:33*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[17*FORCE_DATA_WIDTH-1:16*FORCE_DATA_WIDTH] = force_and_addr[35*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:35*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[17*FORCE_DATA_WIDTH-1:16*FORCE_DATA_WIDTH] = force_and_addr[37*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:37*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[17*FORCE_DATA_WIDTH-1:16*FORCE_DATA_WIDTH] = force_and_addr[44*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:44*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[17*FORCE_DATA_WIDTH-1:16*FORCE_DATA_WIDTH] = force_and_addr[45*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:45*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[17*FORCE_DATA_WIDTH-1:16*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[18*(NUM_NEIGHBOR_CELLS+1)-1:17*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[18*FORCE_DATA_WIDTH-1:17*FORCE_DATA_WIDTH] = force_and_addr[1*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:1*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[18*FORCE_DATA_WIDTH-1:17*FORCE_DATA_WIDTH] = force_and_addr[6*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:6*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[18*FORCE_DATA_WIDTH-1:17*FORCE_DATA_WIDTH] = force_and_addr[13*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:13*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[18*FORCE_DATA_WIDTH-1:17*FORCE_DATA_WIDTH] = force_and_addr[14*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:14*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[18*FORCE_DATA_WIDTH-1:17*FORCE_DATA_WIDTH] = force_and_addr[16*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:16*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[18*FORCE_DATA_WIDTH-1:17*FORCE_DATA_WIDTH] = force_and_addr[17*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:17*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[18*FORCE_DATA_WIDTH-1:17*FORCE_DATA_WIDTH] = force_and_addr[21*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:21*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[18*FORCE_DATA_WIDTH-1:17*FORCE_DATA_WIDTH] = force_and_addr[22*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:22*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[18*FORCE_DATA_WIDTH-1:17*FORCE_DATA_WIDTH] = force_and_addr[30*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:30*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[18*FORCE_DATA_WIDTH-1:17*FORCE_DATA_WIDTH] = force_and_addr[32*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:32*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[18*FORCE_DATA_WIDTH-1:17*FORCE_DATA_WIDTH] = force_and_addr[34*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:34*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[18*FORCE_DATA_WIDTH-1:17*FORCE_DATA_WIDTH] = force_and_addr[38*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:38*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[18*FORCE_DATA_WIDTH-1:17*FORCE_DATA_WIDTH] = force_and_addr[45*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:45*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[18*FORCE_DATA_WIDTH-1:17*FORCE_DATA_WIDTH] = force_and_addr[46*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:46*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[18*FORCE_DATA_WIDTH-1:17*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[19*(NUM_NEIGHBOR_CELLS+1)-1:18*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[19*FORCE_DATA_WIDTH-1:18*FORCE_DATA_WIDTH] = force_and_addr[2*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:2*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[19*FORCE_DATA_WIDTH-1:18*FORCE_DATA_WIDTH] = force_and_addr[7*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:7*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[19*FORCE_DATA_WIDTH-1:18*FORCE_DATA_WIDTH] = force_and_addr[14*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:14*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[19*FORCE_DATA_WIDTH-1:18*FORCE_DATA_WIDTH] = force_and_addr[15*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:15*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[19*FORCE_DATA_WIDTH-1:18*FORCE_DATA_WIDTH] = force_and_addr[17*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:17*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[19*FORCE_DATA_WIDTH-1:18*FORCE_DATA_WIDTH] = force_and_addr[18*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:18*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[19*FORCE_DATA_WIDTH-1:18*FORCE_DATA_WIDTH] = force_and_addr[22*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:22*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[19*FORCE_DATA_WIDTH-1:18*FORCE_DATA_WIDTH] = force_and_addr[23*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:23*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[19*FORCE_DATA_WIDTH-1:18*FORCE_DATA_WIDTH] = force_and_addr[31*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:31*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[19*FORCE_DATA_WIDTH-1:18*FORCE_DATA_WIDTH] = force_and_addr[33*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:33*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[19*FORCE_DATA_WIDTH-1:18*FORCE_DATA_WIDTH] = force_and_addr[35*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:35*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[19*FORCE_DATA_WIDTH-1:18*FORCE_DATA_WIDTH] = force_and_addr[39*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:39*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[19*FORCE_DATA_WIDTH-1:18*FORCE_DATA_WIDTH] = force_and_addr[46*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:46*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[19*FORCE_DATA_WIDTH-1:18*FORCE_DATA_WIDTH] = force_and_addr[47*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:47*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[19*FORCE_DATA_WIDTH-1:18*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[20*(NUM_NEIGHBOR_CELLS+1)-1:19*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[20*FORCE_DATA_WIDTH-1:19*FORCE_DATA_WIDTH] = force_and_addr[3*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:3*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[20*FORCE_DATA_WIDTH-1:19*FORCE_DATA_WIDTH] = force_and_addr[4*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:4*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[20*FORCE_DATA_WIDTH-1:19*FORCE_DATA_WIDTH] = force_and_addr[12*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:12*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[20*FORCE_DATA_WIDTH-1:19*FORCE_DATA_WIDTH] = force_and_addr[15*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:15*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[20*FORCE_DATA_WIDTH-1:19*FORCE_DATA_WIDTH] = force_and_addr[18*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:18*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[20*FORCE_DATA_WIDTH-1:19*FORCE_DATA_WIDTH] = force_and_addr[19*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:19*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[20*FORCE_DATA_WIDTH-1:19*FORCE_DATA_WIDTH] = force_and_addr[20*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:20*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[20*FORCE_DATA_WIDTH-1:19*FORCE_DATA_WIDTH] = force_and_addr[23*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:23*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[20*FORCE_DATA_WIDTH-1:19*FORCE_DATA_WIDTH] = force_and_addr[28*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:28*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[20*FORCE_DATA_WIDTH-1:19*FORCE_DATA_WIDTH] = force_and_addr[32*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:32*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[20*FORCE_DATA_WIDTH-1:19*FORCE_DATA_WIDTH] = force_and_addr[34*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:34*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[20*FORCE_DATA_WIDTH-1:19*FORCE_DATA_WIDTH] = force_and_addr[36*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:36*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[20*FORCE_DATA_WIDTH-1:19*FORCE_DATA_WIDTH] = force_and_addr[44*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:44*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[20*FORCE_DATA_WIDTH-1:19*FORCE_DATA_WIDTH] = force_and_addr[47*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:47*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[20*FORCE_DATA_WIDTH-1:19*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[21*(NUM_NEIGHBOR_CELLS+1)-1:20*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[21*FORCE_DATA_WIDTH-1:20*FORCE_DATA_WIDTH] = force_and_addr[0*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:0*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[21*FORCE_DATA_WIDTH-1:20*FORCE_DATA_WIDTH] = force_and_addr[1*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:1*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[21*FORCE_DATA_WIDTH-1:20*FORCE_DATA_WIDTH] = force_and_addr[4*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:4*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[21*FORCE_DATA_WIDTH-1:20*FORCE_DATA_WIDTH] = force_and_addr[9*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:9*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[21*FORCE_DATA_WIDTH-1:20*FORCE_DATA_WIDTH] = force_and_addr[17*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:17*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[21*FORCE_DATA_WIDTH-1:20*FORCE_DATA_WIDTH] = force_and_addr[20*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:20*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[21*FORCE_DATA_WIDTH-1:20*FORCE_DATA_WIDTH] = force_and_addr[23*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:23*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[21*FORCE_DATA_WIDTH-1:20*FORCE_DATA_WIDTH] = force_and_addr[24*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:24*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[21*FORCE_DATA_WIDTH-1:20*FORCE_DATA_WIDTH] = force_and_addr[25*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:25*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[21*FORCE_DATA_WIDTH-1:20*FORCE_DATA_WIDTH] = force_and_addr[32*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:32*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[21*FORCE_DATA_WIDTH-1:20*FORCE_DATA_WIDTH] = force_and_addr[33*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:33*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[21*FORCE_DATA_WIDTH-1:20*FORCE_DATA_WIDTH] = force_and_addr[37*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:37*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[21*FORCE_DATA_WIDTH-1:20*FORCE_DATA_WIDTH] = force_and_addr[39*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:39*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[21*FORCE_DATA_WIDTH-1:20*FORCE_DATA_WIDTH] = force_and_addr[41*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:41*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[21*FORCE_DATA_WIDTH-1:20*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[22*(NUM_NEIGHBOR_CELLS+1)-1:21*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[22*FORCE_DATA_WIDTH-1:21*FORCE_DATA_WIDTH] = force_and_addr[1*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:1*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[22*FORCE_DATA_WIDTH-1:21*FORCE_DATA_WIDTH] = force_and_addr[2*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:2*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[22*FORCE_DATA_WIDTH-1:21*FORCE_DATA_WIDTH] = force_and_addr[5*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:5*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[22*FORCE_DATA_WIDTH-1:21*FORCE_DATA_WIDTH] = force_and_addr[10*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:10*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[22*FORCE_DATA_WIDTH-1:21*FORCE_DATA_WIDTH] = force_and_addr[18*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:18*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[22*FORCE_DATA_WIDTH-1:21*FORCE_DATA_WIDTH] = force_and_addr[20*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:20*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[22*FORCE_DATA_WIDTH-1:21*FORCE_DATA_WIDTH] = force_and_addr[21*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:21*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[22*FORCE_DATA_WIDTH-1:21*FORCE_DATA_WIDTH] = force_and_addr[25*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:25*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[22*FORCE_DATA_WIDTH-1:21*FORCE_DATA_WIDTH] = force_and_addr[26*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:26*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[22*FORCE_DATA_WIDTH-1:21*FORCE_DATA_WIDTH] = force_and_addr[33*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:33*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[22*FORCE_DATA_WIDTH-1:21*FORCE_DATA_WIDTH] = force_and_addr[34*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:34*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[22*FORCE_DATA_WIDTH-1:21*FORCE_DATA_WIDTH] = force_and_addr[36*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:36*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[22*FORCE_DATA_WIDTH-1:21*FORCE_DATA_WIDTH] = force_and_addr[38*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:38*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[22*FORCE_DATA_WIDTH-1:21*FORCE_DATA_WIDTH] = force_and_addr[42*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:42*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[22*FORCE_DATA_WIDTH-1:21*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[23*(NUM_NEIGHBOR_CELLS+1)-1:22*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[23*FORCE_DATA_WIDTH-1:22*FORCE_DATA_WIDTH] = force_and_addr[2*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:2*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[23*FORCE_DATA_WIDTH-1:22*FORCE_DATA_WIDTH] = force_and_addr[3*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:3*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[23*FORCE_DATA_WIDTH-1:22*FORCE_DATA_WIDTH] = force_and_addr[6*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:6*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[23*FORCE_DATA_WIDTH-1:22*FORCE_DATA_WIDTH] = force_and_addr[11*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:11*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[23*FORCE_DATA_WIDTH-1:22*FORCE_DATA_WIDTH] = force_and_addr[19*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:19*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[23*FORCE_DATA_WIDTH-1:22*FORCE_DATA_WIDTH] = force_and_addr[21*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:21*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[23*FORCE_DATA_WIDTH-1:22*FORCE_DATA_WIDTH] = force_and_addr[22*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:22*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[23*FORCE_DATA_WIDTH-1:22*FORCE_DATA_WIDTH] = force_and_addr[26*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:26*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[23*FORCE_DATA_WIDTH-1:22*FORCE_DATA_WIDTH] = force_and_addr[27*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:27*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[23*FORCE_DATA_WIDTH-1:22*FORCE_DATA_WIDTH] = force_and_addr[34*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:34*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[23*FORCE_DATA_WIDTH-1:22*FORCE_DATA_WIDTH] = force_and_addr[35*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:35*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[23*FORCE_DATA_WIDTH-1:22*FORCE_DATA_WIDTH] = force_and_addr[37*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:37*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[23*FORCE_DATA_WIDTH-1:22*FORCE_DATA_WIDTH] = force_and_addr[39*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:39*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[23*FORCE_DATA_WIDTH-1:22*FORCE_DATA_WIDTH] = force_and_addr[43*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:43*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[23*FORCE_DATA_WIDTH-1:22*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[24*(NUM_NEIGHBOR_CELLS+1)-1:23*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[24*FORCE_DATA_WIDTH-1:23*FORCE_DATA_WIDTH] = force_and_addr[0*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:0*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[24*FORCE_DATA_WIDTH-1:23*FORCE_DATA_WIDTH] = force_and_addr[3*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:3*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[24*FORCE_DATA_WIDTH-1:23*FORCE_DATA_WIDTH] = force_and_addr[7*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:7*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[24*FORCE_DATA_WIDTH-1:23*FORCE_DATA_WIDTH] = force_and_addr[8*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:8*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[24*FORCE_DATA_WIDTH-1:23*FORCE_DATA_WIDTH] = force_and_addr[16*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:16*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[24*FORCE_DATA_WIDTH-1:23*FORCE_DATA_WIDTH] = force_and_addr[22*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:22*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[24*FORCE_DATA_WIDTH-1:23*FORCE_DATA_WIDTH] = force_and_addr[23*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:23*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[24*FORCE_DATA_WIDTH-1:23*FORCE_DATA_WIDTH] = force_and_addr[24*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:24*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[24*FORCE_DATA_WIDTH-1:23*FORCE_DATA_WIDTH] = force_and_addr[27*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:27*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[24*FORCE_DATA_WIDTH-1:23*FORCE_DATA_WIDTH] = force_and_addr[32*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:32*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[24*FORCE_DATA_WIDTH-1:23*FORCE_DATA_WIDTH] = force_and_addr[35*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:35*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[24*FORCE_DATA_WIDTH-1:23*FORCE_DATA_WIDTH] = force_and_addr[36*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:36*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[24*FORCE_DATA_WIDTH-1:23*FORCE_DATA_WIDTH] = force_and_addr[38*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:38*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[24*FORCE_DATA_WIDTH-1:23*FORCE_DATA_WIDTH] = force_and_addr[40*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:40*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[24*FORCE_DATA_WIDTH-1:23*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[25*(NUM_NEIGHBOR_CELLS+1)-1:24*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[25*FORCE_DATA_WIDTH-1:24*FORCE_DATA_WIDTH] = force_and_addr[4*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:4*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[25*FORCE_DATA_WIDTH-1:24*FORCE_DATA_WIDTH] = force_and_addr[5*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:5*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[25*FORCE_DATA_WIDTH-1:24*FORCE_DATA_WIDTH] = force_and_addr[8*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:8*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[25*FORCE_DATA_WIDTH-1:24*FORCE_DATA_WIDTH] = force_and_addr[13*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:13*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[25*FORCE_DATA_WIDTH-1:24*FORCE_DATA_WIDTH] = force_and_addr[21*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:21*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[25*FORCE_DATA_WIDTH-1:24*FORCE_DATA_WIDTH] = force_and_addr[24*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:24*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[25*FORCE_DATA_WIDTH-1:24*FORCE_DATA_WIDTH] = force_and_addr[27*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:27*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[25*FORCE_DATA_WIDTH-1:24*FORCE_DATA_WIDTH] = force_and_addr[28*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:28*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[25*FORCE_DATA_WIDTH-1:24*FORCE_DATA_WIDTH] = force_and_addr[29*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:29*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[25*FORCE_DATA_WIDTH-1:24*FORCE_DATA_WIDTH] = force_and_addr[36*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:36*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[25*FORCE_DATA_WIDTH-1:24*FORCE_DATA_WIDTH] = force_and_addr[37*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:37*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[25*FORCE_DATA_WIDTH-1:24*FORCE_DATA_WIDTH] = force_and_addr[41*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:41*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[25*FORCE_DATA_WIDTH-1:24*FORCE_DATA_WIDTH] = force_and_addr[43*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:43*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[25*FORCE_DATA_WIDTH-1:24*FORCE_DATA_WIDTH] = force_and_addr[45*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:45*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[25*FORCE_DATA_WIDTH-1:24*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[26*(NUM_NEIGHBOR_CELLS+1)-1:25*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[26*FORCE_DATA_WIDTH-1:25*FORCE_DATA_WIDTH] = force_and_addr[5*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:5*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[26*FORCE_DATA_WIDTH-1:25*FORCE_DATA_WIDTH] = force_and_addr[6*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:6*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[26*FORCE_DATA_WIDTH-1:25*FORCE_DATA_WIDTH] = force_and_addr[9*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:9*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[26*FORCE_DATA_WIDTH-1:25*FORCE_DATA_WIDTH] = force_and_addr[14*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:14*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[26*FORCE_DATA_WIDTH-1:25*FORCE_DATA_WIDTH] = force_and_addr[22*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:22*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[26*FORCE_DATA_WIDTH-1:25*FORCE_DATA_WIDTH] = force_and_addr[24*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:24*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[26*FORCE_DATA_WIDTH-1:25*FORCE_DATA_WIDTH] = force_and_addr[25*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:25*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[26*FORCE_DATA_WIDTH-1:25*FORCE_DATA_WIDTH] = force_and_addr[29*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:29*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[26*FORCE_DATA_WIDTH-1:25*FORCE_DATA_WIDTH] = force_and_addr[30*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:30*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[26*FORCE_DATA_WIDTH-1:25*FORCE_DATA_WIDTH] = force_and_addr[37*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:37*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[26*FORCE_DATA_WIDTH-1:25*FORCE_DATA_WIDTH] = force_and_addr[38*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:38*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[26*FORCE_DATA_WIDTH-1:25*FORCE_DATA_WIDTH] = force_and_addr[40*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:40*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[26*FORCE_DATA_WIDTH-1:25*FORCE_DATA_WIDTH] = force_and_addr[42*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:42*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[26*FORCE_DATA_WIDTH-1:25*FORCE_DATA_WIDTH] = force_and_addr[46*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:46*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[26*FORCE_DATA_WIDTH-1:25*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[27*(NUM_NEIGHBOR_CELLS+1)-1:26*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[27*FORCE_DATA_WIDTH-1:26*FORCE_DATA_WIDTH] = force_and_addr[6*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:6*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[27*FORCE_DATA_WIDTH-1:26*FORCE_DATA_WIDTH] = force_and_addr[7*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:7*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[27*FORCE_DATA_WIDTH-1:26*FORCE_DATA_WIDTH] = force_and_addr[10*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:10*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[27*FORCE_DATA_WIDTH-1:26*FORCE_DATA_WIDTH] = force_and_addr[15*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:15*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[27*FORCE_DATA_WIDTH-1:26*FORCE_DATA_WIDTH] = force_and_addr[23*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:23*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[27*FORCE_DATA_WIDTH-1:26*FORCE_DATA_WIDTH] = force_and_addr[25*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:25*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[27*FORCE_DATA_WIDTH-1:26*FORCE_DATA_WIDTH] = force_and_addr[26*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:26*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[27*FORCE_DATA_WIDTH-1:26*FORCE_DATA_WIDTH] = force_and_addr[30*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:30*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[27*FORCE_DATA_WIDTH-1:26*FORCE_DATA_WIDTH] = force_and_addr[31*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:31*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[27*FORCE_DATA_WIDTH-1:26*FORCE_DATA_WIDTH] = force_and_addr[38*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:38*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[27*FORCE_DATA_WIDTH-1:26*FORCE_DATA_WIDTH] = force_and_addr[39*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:39*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[27*FORCE_DATA_WIDTH-1:26*FORCE_DATA_WIDTH] = force_and_addr[41*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:41*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[27*FORCE_DATA_WIDTH-1:26*FORCE_DATA_WIDTH] = force_and_addr[43*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:43*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[27*FORCE_DATA_WIDTH-1:26*FORCE_DATA_WIDTH] = force_and_addr[47*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:47*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[27*FORCE_DATA_WIDTH-1:26*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[28*(NUM_NEIGHBOR_CELLS+1)-1:27*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[28*FORCE_DATA_WIDTH-1:27*FORCE_DATA_WIDTH] = force_and_addr[4*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:4*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[28*FORCE_DATA_WIDTH-1:27*FORCE_DATA_WIDTH] = force_and_addr[7*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:7*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[28*FORCE_DATA_WIDTH-1:27*FORCE_DATA_WIDTH] = force_and_addr[11*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:11*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[28*FORCE_DATA_WIDTH-1:27*FORCE_DATA_WIDTH] = force_and_addr[12*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:12*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[28*FORCE_DATA_WIDTH-1:27*FORCE_DATA_WIDTH] = force_and_addr[20*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:20*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[28*FORCE_DATA_WIDTH-1:27*FORCE_DATA_WIDTH] = force_and_addr[26*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:26*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[28*FORCE_DATA_WIDTH-1:27*FORCE_DATA_WIDTH] = force_and_addr[27*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:27*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[28*FORCE_DATA_WIDTH-1:27*FORCE_DATA_WIDTH] = force_and_addr[28*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:28*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[28*FORCE_DATA_WIDTH-1:27*FORCE_DATA_WIDTH] = force_and_addr[31*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:31*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[28*FORCE_DATA_WIDTH-1:27*FORCE_DATA_WIDTH] = force_and_addr[36*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:36*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[28*FORCE_DATA_WIDTH-1:27*FORCE_DATA_WIDTH] = force_and_addr[39*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:39*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[28*FORCE_DATA_WIDTH-1:27*FORCE_DATA_WIDTH] = force_and_addr[40*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:40*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[28*FORCE_DATA_WIDTH-1:27*FORCE_DATA_WIDTH] = force_and_addr[42*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:42*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[28*FORCE_DATA_WIDTH-1:27*FORCE_DATA_WIDTH] = force_and_addr[44*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:44*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[28*FORCE_DATA_WIDTH-1:27*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[29*(NUM_NEIGHBOR_CELLS+1)-1:28*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[29*FORCE_DATA_WIDTH-1:28*FORCE_DATA_WIDTH] = force_and_addr[1*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:1*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[29*FORCE_DATA_WIDTH-1:28*FORCE_DATA_WIDTH] = force_and_addr[8*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:8*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[29*FORCE_DATA_WIDTH-1:28*FORCE_DATA_WIDTH] = force_and_addr[9*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:9*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[29*FORCE_DATA_WIDTH-1:28*FORCE_DATA_WIDTH] = force_and_addr[12*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:12*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[29*FORCE_DATA_WIDTH-1:28*FORCE_DATA_WIDTH] = force_and_addr[16*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:16*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[29*FORCE_DATA_WIDTH-1:28*FORCE_DATA_WIDTH] = force_and_addr[17*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:17*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[29*FORCE_DATA_WIDTH-1:28*FORCE_DATA_WIDTH] = force_and_addr[25*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:25*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[29*FORCE_DATA_WIDTH-1:28*FORCE_DATA_WIDTH] = force_and_addr[28*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:28*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[29*FORCE_DATA_WIDTH-1:28*FORCE_DATA_WIDTH] = force_and_addr[31*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:31*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[29*FORCE_DATA_WIDTH-1:28*FORCE_DATA_WIDTH] = force_and_addr[33*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:33*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[29*FORCE_DATA_WIDTH-1:28*FORCE_DATA_WIDTH] = force_and_addr[40*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:40*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[29*FORCE_DATA_WIDTH-1:28*FORCE_DATA_WIDTH] = force_and_addr[41*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:41*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[29*FORCE_DATA_WIDTH-1:28*FORCE_DATA_WIDTH] = force_and_addr[45*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:45*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[29*FORCE_DATA_WIDTH-1:28*FORCE_DATA_WIDTH] = force_and_addr[47*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:47*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[29*FORCE_DATA_WIDTH-1:28*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[30*(NUM_NEIGHBOR_CELLS+1)-1:29*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[30*FORCE_DATA_WIDTH-1:29*FORCE_DATA_WIDTH] = force_and_addr[2*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:2*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[30*FORCE_DATA_WIDTH-1:29*FORCE_DATA_WIDTH] = force_and_addr[9*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:9*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[30*FORCE_DATA_WIDTH-1:29*FORCE_DATA_WIDTH] = force_and_addr[10*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:10*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[30*FORCE_DATA_WIDTH-1:29*FORCE_DATA_WIDTH] = force_and_addr[13*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:13*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[30*FORCE_DATA_WIDTH-1:29*FORCE_DATA_WIDTH] = force_and_addr[17*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:17*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[30*FORCE_DATA_WIDTH-1:29*FORCE_DATA_WIDTH] = force_and_addr[18*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:18*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[30*FORCE_DATA_WIDTH-1:29*FORCE_DATA_WIDTH] = force_and_addr[26*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:26*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[30*FORCE_DATA_WIDTH-1:29*FORCE_DATA_WIDTH] = force_and_addr[28*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:28*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[30*FORCE_DATA_WIDTH-1:29*FORCE_DATA_WIDTH] = force_and_addr[29*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:29*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[30*FORCE_DATA_WIDTH-1:29*FORCE_DATA_WIDTH] = force_and_addr[34*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:34*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[30*FORCE_DATA_WIDTH-1:29*FORCE_DATA_WIDTH] = force_and_addr[41*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:41*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[30*FORCE_DATA_WIDTH-1:29*FORCE_DATA_WIDTH] = force_and_addr[42*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:42*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[30*FORCE_DATA_WIDTH-1:29*FORCE_DATA_WIDTH] = force_and_addr[44*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:44*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[30*FORCE_DATA_WIDTH-1:29*FORCE_DATA_WIDTH] = force_and_addr[46*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:46*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[30*FORCE_DATA_WIDTH-1:29*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[31*(NUM_NEIGHBOR_CELLS+1)-1:30*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[31*FORCE_DATA_WIDTH-1:30*FORCE_DATA_WIDTH] = force_and_addr[3*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:3*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[31*FORCE_DATA_WIDTH-1:30*FORCE_DATA_WIDTH] = force_and_addr[10*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:10*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[31*FORCE_DATA_WIDTH-1:30*FORCE_DATA_WIDTH] = force_and_addr[11*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:11*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[31*FORCE_DATA_WIDTH-1:30*FORCE_DATA_WIDTH] = force_and_addr[14*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:14*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[31*FORCE_DATA_WIDTH-1:30*FORCE_DATA_WIDTH] = force_and_addr[18*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:18*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[31*FORCE_DATA_WIDTH-1:30*FORCE_DATA_WIDTH] = force_and_addr[19*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:19*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[31*FORCE_DATA_WIDTH-1:30*FORCE_DATA_WIDTH] = force_and_addr[27*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:27*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[31*FORCE_DATA_WIDTH-1:30*FORCE_DATA_WIDTH] = force_and_addr[29*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:29*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[31*FORCE_DATA_WIDTH-1:30*FORCE_DATA_WIDTH] = force_and_addr[30*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:30*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[31*FORCE_DATA_WIDTH-1:30*FORCE_DATA_WIDTH] = force_and_addr[35*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:35*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[31*FORCE_DATA_WIDTH-1:30*FORCE_DATA_WIDTH] = force_and_addr[42*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:42*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[31*FORCE_DATA_WIDTH-1:30*FORCE_DATA_WIDTH] = force_and_addr[43*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:43*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[31*FORCE_DATA_WIDTH-1:30*FORCE_DATA_WIDTH] = force_and_addr[45*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:45*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[31*FORCE_DATA_WIDTH-1:30*FORCE_DATA_WIDTH] = force_and_addr[47*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:47*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[31*FORCE_DATA_WIDTH-1:30*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[32*(NUM_NEIGHBOR_CELLS+1)-1:31*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[32*FORCE_DATA_WIDTH-1:31*FORCE_DATA_WIDTH] = force_and_addr[0*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:0*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[32*FORCE_DATA_WIDTH-1:31*FORCE_DATA_WIDTH] = force_and_addr[8*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:8*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[32*FORCE_DATA_WIDTH-1:31*FORCE_DATA_WIDTH] = force_and_addr[11*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:11*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[32*FORCE_DATA_WIDTH-1:31*FORCE_DATA_WIDTH] = force_and_addr[15*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:15*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[32*FORCE_DATA_WIDTH-1:31*FORCE_DATA_WIDTH] = force_and_addr[16*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:16*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[32*FORCE_DATA_WIDTH-1:31*FORCE_DATA_WIDTH] = force_and_addr[19*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:19*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[32*FORCE_DATA_WIDTH-1:31*FORCE_DATA_WIDTH] = force_and_addr[24*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:24*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[32*FORCE_DATA_WIDTH-1:31*FORCE_DATA_WIDTH] = force_and_addr[30*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:30*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[32*FORCE_DATA_WIDTH-1:31*FORCE_DATA_WIDTH] = force_and_addr[31*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:31*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[32*FORCE_DATA_WIDTH-1:31*FORCE_DATA_WIDTH] = force_and_addr[32*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:32*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[32*FORCE_DATA_WIDTH-1:31*FORCE_DATA_WIDTH] = force_and_addr[40*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:40*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[32*FORCE_DATA_WIDTH-1:31*FORCE_DATA_WIDTH] = force_and_addr[43*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:43*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[32*FORCE_DATA_WIDTH-1:31*FORCE_DATA_WIDTH] = force_and_addr[44*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:44*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[32*FORCE_DATA_WIDTH-1:31*FORCE_DATA_WIDTH] = force_and_addr[46*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:46*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[32*FORCE_DATA_WIDTH-1:31*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[33*(NUM_NEIGHBOR_CELLS+1)-1:32*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[33*FORCE_DATA_WIDTH-1:32*FORCE_DATA_WIDTH] = force_and_addr[16*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:16*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[33*FORCE_DATA_WIDTH-1:32*FORCE_DATA_WIDTH] = force_and_addr[21*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:21*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[33*FORCE_DATA_WIDTH-1:32*FORCE_DATA_WIDTH] = force_and_addr[28*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:28*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[33*FORCE_DATA_WIDTH-1:32*FORCE_DATA_WIDTH] = force_and_addr[29*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:29*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[33*FORCE_DATA_WIDTH-1:32*FORCE_DATA_WIDTH] = force_and_addr[32*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:32*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[33*FORCE_DATA_WIDTH-1:32*FORCE_DATA_WIDTH] = force_and_addr[35*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:35*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[33*FORCE_DATA_WIDTH-1:32*FORCE_DATA_WIDTH] = force_and_addr[36*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:36*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[33*FORCE_DATA_WIDTH-1:32*FORCE_DATA_WIDTH] = force_and_addr[37*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:37*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[33*FORCE_DATA_WIDTH-1:32*FORCE_DATA_WIDTH] = force_and_addr[45*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:45*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[33*FORCE_DATA_WIDTH-1:32*FORCE_DATA_WIDTH] = force_and_addr[49*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:49*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[33*FORCE_DATA_WIDTH-1:32*FORCE_DATA_WIDTH] = force_and_addr[51*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:51*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[33*FORCE_DATA_WIDTH-1:32*FORCE_DATA_WIDTH] = force_and_addr[53*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:53*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[33*FORCE_DATA_WIDTH-1:32*FORCE_DATA_WIDTH] = force_and_addr[60*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:60*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[33*FORCE_DATA_WIDTH-1:32*FORCE_DATA_WIDTH] = force_and_addr[61*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:61*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[33*FORCE_DATA_WIDTH-1:32*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[34*(NUM_NEIGHBOR_CELLS+1)-1:33*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[34*FORCE_DATA_WIDTH-1:33*FORCE_DATA_WIDTH] = force_and_addr[17*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:17*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[34*FORCE_DATA_WIDTH-1:33*FORCE_DATA_WIDTH] = force_and_addr[22*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:22*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[34*FORCE_DATA_WIDTH-1:33*FORCE_DATA_WIDTH] = force_and_addr[29*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:29*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[34*FORCE_DATA_WIDTH-1:33*FORCE_DATA_WIDTH] = force_and_addr[30*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:30*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[34*FORCE_DATA_WIDTH-1:33*FORCE_DATA_WIDTH] = force_and_addr[32*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:32*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[34*FORCE_DATA_WIDTH-1:33*FORCE_DATA_WIDTH] = force_and_addr[33*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:33*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[34*FORCE_DATA_WIDTH-1:33*FORCE_DATA_WIDTH] = force_and_addr[37*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:37*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[34*FORCE_DATA_WIDTH-1:33*FORCE_DATA_WIDTH] = force_and_addr[38*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:38*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[34*FORCE_DATA_WIDTH-1:33*FORCE_DATA_WIDTH] = force_and_addr[46*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:46*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[34*FORCE_DATA_WIDTH-1:33*FORCE_DATA_WIDTH] = force_and_addr[48*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:48*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[34*FORCE_DATA_WIDTH-1:33*FORCE_DATA_WIDTH] = force_and_addr[50*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:50*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[34*FORCE_DATA_WIDTH-1:33*FORCE_DATA_WIDTH] = force_and_addr[54*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:54*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[34*FORCE_DATA_WIDTH-1:33*FORCE_DATA_WIDTH] = force_and_addr[61*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:61*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[34*FORCE_DATA_WIDTH-1:33*FORCE_DATA_WIDTH] = force_and_addr[62*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:62*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[34*FORCE_DATA_WIDTH-1:33*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[35*(NUM_NEIGHBOR_CELLS+1)-1:34*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[35*FORCE_DATA_WIDTH-1:34*FORCE_DATA_WIDTH] = force_and_addr[18*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:18*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[35*FORCE_DATA_WIDTH-1:34*FORCE_DATA_WIDTH] = force_and_addr[23*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:23*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[35*FORCE_DATA_WIDTH-1:34*FORCE_DATA_WIDTH] = force_and_addr[30*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:30*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[35*FORCE_DATA_WIDTH-1:34*FORCE_DATA_WIDTH] = force_and_addr[31*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:31*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[35*FORCE_DATA_WIDTH-1:34*FORCE_DATA_WIDTH] = force_and_addr[33*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:33*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[35*FORCE_DATA_WIDTH-1:34*FORCE_DATA_WIDTH] = force_and_addr[34*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:34*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[35*FORCE_DATA_WIDTH-1:34*FORCE_DATA_WIDTH] = force_and_addr[38*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:38*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[35*FORCE_DATA_WIDTH-1:34*FORCE_DATA_WIDTH] = force_and_addr[39*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:39*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[35*FORCE_DATA_WIDTH-1:34*FORCE_DATA_WIDTH] = force_and_addr[47*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:47*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[35*FORCE_DATA_WIDTH-1:34*FORCE_DATA_WIDTH] = force_and_addr[49*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:49*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[35*FORCE_DATA_WIDTH-1:34*FORCE_DATA_WIDTH] = force_and_addr[51*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:51*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[35*FORCE_DATA_WIDTH-1:34*FORCE_DATA_WIDTH] = force_and_addr[55*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:55*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[35*FORCE_DATA_WIDTH-1:34*FORCE_DATA_WIDTH] = force_and_addr[62*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:62*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[35*FORCE_DATA_WIDTH-1:34*FORCE_DATA_WIDTH] = force_and_addr[63*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:63*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[35*FORCE_DATA_WIDTH-1:34*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[36*(NUM_NEIGHBOR_CELLS+1)-1:35*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[36*FORCE_DATA_WIDTH-1:35*FORCE_DATA_WIDTH] = force_and_addr[19*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:19*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[36*FORCE_DATA_WIDTH-1:35*FORCE_DATA_WIDTH] = force_and_addr[20*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:20*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[36*FORCE_DATA_WIDTH-1:35*FORCE_DATA_WIDTH] = force_and_addr[28*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:28*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[36*FORCE_DATA_WIDTH-1:35*FORCE_DATA_WIDTH] = force_and_addr[31*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:31*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[36*FORCE_DATA_WIDTH-1:35*FORCE_DATA_WIDTH] = force_and_addr[34*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:34*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[36*FORCE_DATA_WIDTH-1:35*FORCE_DATA_WIDTH] = force_and_addr[35*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:35*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[36*FORCE_DATA_WIDTH-1:35*FORCE_DATA_WIDTH] = force_and_addr[36*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:36*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[36*FORCE_DATA_WIDTH-1:35*FORCE_DATA_WIDTH] = force_and_addr[39*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:39*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[36*FORCE_DATA_WIDTH-1:35*FORCE_DATA_WIDTH] = force_and_addr[44*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:44*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[36*FORCE_DATA_WIDTH-1:35*FORCE_DATA_WIDTH] = force_and_addr[48*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:48*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[36*FORCE_DATA_WIDTH-1:35*FORCE_DATA_WIDTH] = force_and_addr[50*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:50*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[36*FORCE_DATA_WIDTH-1:35*FORCE_DATA_WIDTH] = force_and_addr[52*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:52*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[36*FORCE_DATA_WIDTH-1:35*FORCE_DATA_WIDTH] = force_and_addr[60*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:60*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[36*FORCE_DATA_WIDTH-1:35*FORCE_DATA_WIDTH] = force_and_addr[63*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:63*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[36*FORCE_DATA_WIDTH-1:35*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[37*(NUM_NEIGHBOR_CELLS+1)-1:36*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[37*FORCE_DATA_WIDTH-1:36*FORCE_DATA_WIDTH] = force_and_addr[16*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:16*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[37*FORCE_DATA_WIDTH-1:36*FORCE_DATA_WIDTH] = force_and_addr[17*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:17*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[37*FORCE_DATA_WIDTH-1:36*FORCE_DATA_WIDTH] = force_and_addr[20*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:20*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[37*FORCE_DATA_WIDTH-1:36*FORCE_DATA_WIDTH] = force_and_addr[25*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:25*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[37*FORCE_DATA_WIDTH-1:36*FORCE_DATA_WIDTH] = force_and_addr[33*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:33*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[37*FORCE_DATA_WIDTH-1:36*FORCE_DATA_WIDTH] = force_and_addr[36*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:36*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[37*FORCE_DATA_WIDTH-1:36*FORCE_DATA_WIDTH] = force_and_addr[39*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:39*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[37*FORCE_DATA_WIDTH-1:36*FORCE_DATA_WIDTH] = force_and_addr[40*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:40*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[37*FORCE_DATA_WIDTH-1:36*FORCE_DATA_WIDTH] = force_and_addr[41*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:41*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[37*FORCE_DATA_WIDTH-1:36*FORCE_DATA_WIDTH] = force_and_addr[48*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:48*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[37*FORCE_DATA_WIDTH-1:36*FORCE_DATA_WIDTH] = force_and_addr[49*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:49*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[37*FORCE_DATA_WIDTH-1:36*FORCE_DATA_WIDTH] = force_and_addr[53*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:53*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[37*FORCE_DATA_WIDTH-1:36*FORCE_DATA_WIDTH] = force_and_addr[55*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:55*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[37*FORCE_DATA_WIDTH-1:36*FORCE_DATA_WIDTH] = force_and_addr[57*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:57*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[37*FORCE_DATA_WIDTH-1:36*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[38*(NUM_NEIGHBOR_CELLS+1)-1:37*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[38*FORCE_DATA_WIDTH-1:37*FORCE_DATA_WIDTH] = force_and_addr[17*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:17*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[38*FORCE_DATA_WIDTH-1:37*FORCE_DATA_WIDTH] = force_and_addr[18*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:18*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[38*FORCE_DATA_WIDTH-1:37*FORCE_DATA_WIDTH] = force_and_addr[21*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:21*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[38*FORCE_DATA_WIDTH-1:37*FORCE_DATA_WIDTH] = force_and_addr[26*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:26*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[38*FORCE_DATA_WIDTH-1:37*FORCE_DATA_WIDTH] = force_and_addr[34*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:34*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[38*FORCE_DATA_WIDTH-1:37*FORCE_DATA_WIDTH] = force_and_addr[36*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:36*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[38*FORCE_DATA_WIDTH-1:37*FORCE_DATA_WIDTH] = force_and_addr[37*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:37*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[38*FORCE_DATA_WIDTH-1:37*FORCE_DATA_WIDTH] = force_and_addr[41*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:41*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[38*FORCE_DATA_WIDTH-1:37*FORCE_DATA_WIDTH] = force_and_addr[42*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:42*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[38*FORCE_DATA_WIDTH-1:37*FORCE_DATA_WIDTH] = force_and_addr[49*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:49*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[38*FORCE_DATA_WIDTH-1:37*FORCE_DATA_WIDTH] = force_and_addr[50*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:50*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[38*FORCE_DATA_WIDTH-1:37*FORCE_DATA_WIDTH] = force_and_addr[52*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:52*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[38*FORCE_DATA_WIDTH-1:37*FORCE_DATA_WIDTH] = force_and_addr[54*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:54*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[38*FORCE_DATA_WIDTH-1:37*FORCE_DATA_WIDTH] = force_and_addr[58*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:58*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[38*FORCE_DATA_WIDTH-1:37*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[39*(NUM_NEIGHBOR_CELLS+1)-1:38*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[39*FORCE_DATA_WIDTH-1:38*FORCE_DATA_WIDTH] = force_and_addr[18*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:18*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[39*FORCE_DATA_WIDTH-1:38*FORCE_DATA_WIDTH] = force_and_addr[19*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:19*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[39*FORCE_DATA_WIDTH-1:38*FORCE_DATA_WIDTH] = force_and_addr[22*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:22*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[39*FORCE_DATA_WIDTH-1:38*FORCE_DATA_WIDTH] = force_and_addr[27*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:27*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[39*FORCE_DATA_WIDTH-1:38*FORCE_DATA_WIDTH] = force_and_addr[35*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:35*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[39*FORCE_DATA_WIDTH-1:38*FORCE_DATA_WIDTH] = force_and_addr[37*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:37*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[39*FORCE_DATA_WIDTH-1:38*FORCE_DATA_WIDTH] = force_and_addr[38*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:38*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[39*FORCE_DATA_WIDTH-1:38*FORCE_DATA_WIDTH] = force_and_addr[42*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:42*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[39*FORCE_DATA_WIDTH-1:38*FORCE_DATA_WIDTH] = force_and_addr[43*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:43*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[39*FORCE_DATA_WIDTH-1:38*FORCE_DATA_WIDTH] = force_and_addr[50*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:50*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[39*FORCE_DATA_WIDTH-1:38*FORCE_DATA_WIDTH] = force_and_addr[51*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:51*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[39*FORCE_DATA_WIDTH-1:38*FORCE_DATA_WIDTH] = force_and_addr[53*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:53*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[39*FORCE_DATA_WIDTH-1:38*FORCE_DATA_WIDTH] = force_and_addr[55*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:55*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[39*FORCE_DATA_WIDTH-1:38*FORCE_DATA_WIDTH] = force_and_addr[59*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:59*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[39*FORCE_DATA_WIDTH-1:38*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[40*(NUM_NEIGHBOR_CELLS+1)-1:39*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[40*FORCE_DATA_WIDTH-1:39*FORCE_DATA_WIDTH] = force_and_addr[16*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:16*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[40*FORCE_DATA_WIDTH-1:39*FORCE_DATA_WIDTH] = force_and_addr[19*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:19*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[40*FORCE_DATA_WIDTH-1:39*FORCE_DATA_WIDTH] = force_and_addr[23*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:23*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[40*FORCE_DATA_WIDTH-1:39*FORCE_DATA_WIDTH] = force_and_addr[24*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:24*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[40*FORCE_DATA_WIDTH-1:39*FORCE_DATA_WIDTH] = force_and_addr[32*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:32*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[40*FORCE_DATA_WIDTH-1:39*FORCE_DATA_WIDTH] = force_and_addr[38*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:38*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[40*FORCE_DATA_WIDTH-1:39*FORCE_DATA_WIDTH] = force_and_addr[39*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:39*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[40*FORCE_DATA_WIDTH-1:39*FORCE_DATA_WIDTH] = force_and_addr[40*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:40*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[40*FORCE_DATA_WIDTH-1:39*FORCE_DATA_WIDTH] = force_and_addr[43*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:43*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[40*FORCE_DATA_WIDTH-1:39*FORCE_DATA_WIDTH] = force_and_addr[48*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:48*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[40*FORCE_DATA_WIDTH-1:39*FORCE_DATA_WIDTH] = force_and_addr[51*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:51*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[40*FORCE_DATA_WIDTH-1:39*FORCE_DATA_WIDTH] = force_and_addr[52*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:52*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[40*FORCE_DATA_WIDTH-1:39*FORCE_DATA_WIDTH] = force_and_addr[54*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:54*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[40*FORCE_DATA_WIDTH-1:39*FORCE_DATA_WIDTH] = force_and_addr[56*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:56*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[40*FORCE_DATA_WIDTH-1:39*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[41*(NUM_NEIGHBOR_CELLS+1)-1:40*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[41*FORCE_DATA_WIDTH-1:40*FORCE_DATA_WIDTH] = force_and_addr[20*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:20*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[41*FORCE_DATA_WIDTH-1:40*FORCE_DATA_WIDTH] = force_and_addr[21*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:21*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[41*FORCE_DATA_WIDTH-1:40*FORCE_DATA_WIDTH] = force_and_addr[24*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:24*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[41*FORCE_DATA_WIDTH-1:40*FORCE_DATA_WIDTH] = force_and_addr[29*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:29*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[41*FORCE_DATA_WIDTH-1:40*FORCE_DATA_WIDTH] = force_and_addr[37*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:37*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[41*FORCE_DATA_WIDTH-1:40*FORCE_DATA_WIDTH] = force_and_addr[40*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:40*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[41*FORCE_DATA_WIDTH-1:40*FORCE_DATA_WIDTH] = force_and_addr[43*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:43*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[41*FORCE_DATA_WIDTH-1:40*FORCE_DATA_WIDTH] = force_and_addr[44*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:44*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[41*FORCE_DATA_WIDTH-1:40*FORCE_DATA_WIDTH] = force_and_addr[45*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:45*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[41*FORCE_DATA_WIDTH-1:40*FORCE_DATA_WIDTH] = force_and_addr[52*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:52*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[41*FORCE_DATA_WIDTH-1:40*FORCE_DATA_WIDTH] = force_and_addr[53*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:53*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[41*FORCE_DATA_WIDTH-1:40*FORCE_DATA_WIDTH] = force_and_addr[57*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:57*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[41*FORCE_DATA_WIDTH-1:40*FORCE_DATA_WIDTH] = force_and_addr[59*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:59*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[41*FORCE_DATA_WIDTH-1:40*FORCE_DATA_WIDTH] = force_and_addr[61*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:61*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[41*FORCE_DATA_WIDTH-1:40*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[42*(NUM_NEIGHBOR_CELLS+1)-1:41*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[42*FORCE_DATA_WIDTH-1:41*FORCE_DATA_WIDTH] = force_and_addr[21*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:21*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[42*FORCE_DATA_WIDTH-1:41*FORCE_DATA_WIDTH] = force_and_addr[22*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:22*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[42*FORCE_DATA_WIDTH-1:41*FORCE_DATA_WIDTH] = force_and_addr[25*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:25*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[42*FORCE_DATA_WIDTH-1:41*FORCE_DATA_WIDTH] = force_and_addr[30*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:30*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[42*FORCE_DATA_WIDTH-1:41*FORCE_DATA_WIDTH] = force_and_addr[38*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:38*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[42*FORCE_DATA_WIDTH-1:41*FORCE_DATA_WIDTH] = force_and_addr[40*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:40*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[42*FORCE_DATA_WIDTH-1:41*FORCE_DATA_WIDTH] = force_and_addr[41*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:41*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[42*FORCE_DATA_WIDTH-1:41*FORCE_DATA_WIDTH] = force_and_addr[45*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:45*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[42*FORCE_DATA_WIDTH-1:41*FORCE_DATA_WIDTH] = force_and_addr[46*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:46*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[42*FORCE_DATA_WIDTH-1:41*FORCE_DATA_WIDTH] = force_and_addr[53*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:53*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[42*FORCE_DATA_WIDTH-1:41*FORCE_DATA_WIDTH] = force_and_addr[54*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:54*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[42*FORCE_DATA_WIDTH-1:41*FORCE_DATA_WIDTH] = force_and_addr[56*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:56*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[42*FORCE_DATA_WIDTH-1:41*FORCE_DATA_WIDTH] = force_and_addr[58*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:58*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[42*FORCE_DATA_WIDTH-1:41*FORCE_DATA_WIDTH] = force_and_addr[62*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:62*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[42*FORCE_DATA_WIDTH-1:41*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[43*(NUM_NEIGHBOR_CELLS+1)-1:42*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[43*FORCE_DATA_WIDTH-1:42*FORCE_DATA_WIDTH] = force_and_addr[22*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:22*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[43*FORCE_DATA_WIDTH-1:42*FORCE_DATA_WIDTH] = force_and_addr[23*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:23*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[43*FORCE_DATA_WIDTH-1:42*FORCE_DATA_WIDTH] = force_and_addr[26*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:26*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[43*FORCE_DATA_WIDTH-1:42*FORCE_DATA_WIDTH] = force_and_addr[31*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:31*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[43*FORCE_DATA_WIDTH-1:42*FORCE_DATA_WIDTH] = force_and_addr[39*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:39*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[43*FORCE_DATA_WIDTH-1:42*FORCE_DATA_WIDTH] = force_and_addr[41*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:41*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[43*FORCE_DATA_WIDTH-1:42*FORCE_DATA_WIDTH] = force_and_addr[42*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:42*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[43*FORCE_DATA_WIDTH-1:42*FORCE_DATA_WIDTH] = force_and_addr[46*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:46*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[43*FORCE_DATA_WIDTH-1:42*FORCE_DATA_WIDTH] = force_and_addr[47*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:47*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[43*FORCE_DATA_WIDTH-1:42*FORCE_DATA_WIDTH] = force_and_addr[54*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:54*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[43*FORCE_DATA_WIDTH-1:42*FORCE_DATA_WIDTH] = force_and_addr[55*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:55*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[43*FORCE_DATA_WIDTH-1:42*FORCE_DATA_WIDTH] = force_and_addr[57*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:57*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[43*FORCE_DATA_WIDTH-1:42*FORCE_DATA_WIDTH] = force_and_addr[59*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:59*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[43*FORCE_DATA_WIDTH-1:42*FORCE_DATA_WIDTH] = force_and_addr[63*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:63*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[43*FORCE_DATA_WIDTH-1:42*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[44*(NUM_NEIGHBOR_CELLS+1)-1:43*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[44*FORCE_DATA_WIDTH-1:43*FORCE_DATA_WIDTH] = force_and_addr[20*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:20*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[44*FORCE_DATA_WIDTH-1:43*FORCE_DATA_WIDTH] = force_and_addr[23*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:23*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[44*FORCE_DATA_WIDTH-1:43*FORCE_DATA_WIDTH] = force_and_addr[27*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:27*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[44*FORCE_DATA_WIDTH-1:43*FORCE_DATA_WIDTH] = force_and_addr[28*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:28*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[44*FORCE_DATA_WIDTH-1:43*FORCE_DATA_WIDTH] = force_and_addr[36*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:36*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[44*FORCE_DATA_WIDTH-1:43*FORCE_DATA_WIDTH] = force_and_addr[42*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:42*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[44*FORCE_DATA_WIDTH-1:43*FORCE_DATA_WIDTH] = force_and_addr[43*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:43*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[44*FORCE_DATA_WIDTH-1:43*FORCE_DATA_WIDTH] = force_and_addr[44*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:44*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[44*FORCE_DATA_WIDTH-1:43*FORCE_DATA_WIDTH] = force_and_addr[47*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:47*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[44*FORCE_DATA_WIDTH-1:43*FORCE_DATA_WIDTH] = force_and_addr[52*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:52*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[44*FORCE_DATA_WIDTH-1:43*FORCE_DATA_WIDTH] = force_and_addr[55*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:55*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[44*FORCE_DATA_WIDTH-1:43*FORCE_DATA_WIDTH] = force_and_addr[56*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:56*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[44*FORCE_DATA_WIDTH-1:43*FORCE_DATA_WIDTH] = force_and_addr[58*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:58*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[44*FORCE_DATA_WIDTH-1:43*FORCE_DATA_WIDTH] = force_and_addr[60*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:60*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[44*FORCE_DATA_WIDTH-1:43*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[45*(NUM_NEIGHBOR_CELLS+1)-1:44*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[45*FORCE_DATA_WIDTH-1:44*FORCE_DATA_WIDTH] = force_and_addr[17*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:17*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[45*FORCE_DATA_WIDTH-1:44*FORCE_DATA_WIDTH] = force_and_addr[24*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:24*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[45*FORCE_DATA_WIDTH-1:44*FORCE_DATA_WIDTH] = force_and_addr[25*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:25*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[45*FORCE_DATA_WIDTH-1:44*FORCE_DATA_WIDTH] = force_and_addr[28*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:28*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[45*FORCE_DATA_WIDTH-1:44*FORCE_DATA_WIDTH] = force_and_addr[32*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:32*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[45*FORCE_DATA_WIDTH-1:44*FORCE_DATA_WIDTH] = force_and_addr[33*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:33*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[45*FORCE_DATA_WIDTH-1:44*FORCE_DATA_WIDTH] = force_and_addr[41*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:41*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[45*FORCE_DATA_WIDTH-1:44*FORCE_DATA_WIDTH] = force_and_addr[44*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:44*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[45*FORCE_DATA_WIDTH-1:44*FORCE_DATA_WIDTH] = force_and_addr[47*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:47*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[45*FORCE_DATA_WIDTH-1:44*FORCE_DATA_WIDTH] = force_and_addr[49*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:49*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[45*FORCE_DATA_WIDTH-1:44*FORCE_DATA_WIDTH] = force_and_addr[56*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:56*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[45*FORCE_DATA_WIDTH-1:44*FORCE_DATA_WIDTH] = force_and_addr[57*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:57*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[45*FORCE_DATA_WIDTH-1:44*FORCE_DATA_WIDTH] = force_and_addr[61*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:61*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[45*FORCE_DATA_WIDTH-1:44*FORCE_DATA_WIDTH] = force_and_addr[63*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:63*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[45*FORCE_DATA_WIDTH-1:44*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[46*(NUM_NEIGHBOR_CELLS+1)-1:45*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[46*FORCE_DATA_WIDTH-1:45*FORCE_DATA_WIDTH] = force_and_addr[18*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:18*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[46*FORCE_DATA_WIDTH-1:45*FORCE_DATA_WIDTH] = force_and_addr[25*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:25*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[46*FORCE_DATA_WIDTH-1:45*FORCE_DATA_WIDTH] = force_and_addr[26*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:26*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[46*FORCE_DATA_WIDTH-1:45*FORCE_DATA_WIDTH] = force_and_addr[29*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:29*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[46*FORCE_DATA_WIDTH-1:45*FORCE_DATA_WIDTH] = force_and_addr[33*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:33*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[46*FORCE_DATA_WIDTH-1:45*FORCE_DATA_WIDTH] = force_and_addr[34*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:34*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[46*FORCE_DATA_WIDTH-1:45*FORCE_DATA_WIDTH] = force_and_addr[42*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:42*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[46*FORCE_DATA_WIDTH-1:45*FORCE_DATA_WIDTH] = force_and_addr[44*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:44*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[46*FORCE_DATA_WIDTH-1:45*FORCE_DATA_WIDTH] = force_and_addr[45*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:45*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[46*FORCE_DATA_WIDTH-1:45*FORCE_DATA_WIDTH] = force_and_addr[50*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:50*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[46*FORCE_DATA_WIDTH-1:45*FORCE_DATA_WIDTH] = force_and_addr[57*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:57*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[46*FORCE_DATA_WIDTH-1:45*FORCE_DATA_WIDTH] = force_and_addr[58*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:58*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[46*FORCE_DATA_WIDTH-1:45*FORCE_DATA_WIDTH] = force_and_addr[60*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:60*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[46*FORCE_DATA_WIDTH-1:45*FORCE_DATA_WIDTH] = force_and_addr[62*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:62*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[46*FORCE_DATA_WIDTH-1:45*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[47*(NUM_NEIGHBOR_CELLS+1)-1:46*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[47*FORCE_DATA_WIDTH-1:46*FORCE_DATA_WIDTH] = force_and_addr[19*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:19*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[47*FORCE_DATA_WIDTH-1:46*FORCE_DATA_WIDTH] = force_and_addr[26*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:26*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[47*FORCE_DATA_WIDTH-1:46*FORCE_DATA_WIDTH] = force_and_addr[27*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:27*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[47*FORCE_DATA_WIDTH-1:46*FORCE_DATA_WIDTH] = force_and_addr[30*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:30*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[47*FORCE_DATA_WIDTH-1:46*FORCE_DATA_WIDTH] = force_and_addr[34*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:34*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[47*FORCE_DATA_WIDTH-1:46*FORCE_DATA_WIDTH] = force_and_addr[35*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:35*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[47*FORCE_DATA_WIDTH-1:46*FORCE_DATA_WIDTH] = force_and_addr[43*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:43*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[47*FORCE_DATA_WIDTH-1:46*FORCE_DATA_WIDTH] = force_and_addr[45*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:45*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[47*FORCE_DATA_WIDTH-1:46*FORCE_DATA_WIDTH] = force_and_addr[46*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:46*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[47*FORCE_DATA_WIDTH-1:46*FORCE_DATA_WIDTH] = force_and_addr[51*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:51*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[47*FORCE_DATA_WIDTH-1:46*FORCE_DATA_WIDTH] = force_and_addr[58*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:58*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[47*FORCE_DATA_WIDTH-1:46*FORCE_DATA_WIDTH] = force_and_addr[59*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:59*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[47*FORCE_DATA_WIDTH-1:46*FORCE_DATA_WIDTH] = force_and_addr[61*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:61*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[47*FORCE_DATA_WIDTH-1:46*FORCE_DATA_WIDTH] = force_and_addr[63*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:63*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[47*FORCE_DATA_WIDTH-1:46*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[48*(NUM_NEIGHBOR_CELLS+1)-1:47*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[48*FORCE_DATA_WIDTH-1:47*FORCE_DATA_WIDTH] = force_and_addr[16*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:16*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[48*FORCE_DATA_WIDTH-1:47*FORCE_DATA_WIDTH] = force_and_addr[24*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:24*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[48*FORCE_DATA_WIDTH-1:47*FORCE_DATA_WIDTH] = force_and_addr[27*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:27*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[48*FORCE_DATA_WIDTH-1:47*FORCE_DATA_WIDTH] = force_and_addr[31*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:31*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[48*FORCE_DATA_WIDTH-1:47*FORCE_DATA_WIDTH] = force_and_addr[32*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:32*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[48*FORCE_DATA_WIDTH-1:47*FORCE_DATA_WIDTH] = force_and_addr[35*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:35*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[48*FORCE_DATA_WIDTH-1:47*FORCE_DATA_WIDTH] = force_and_addr[40*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:40*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[48*FORCE_DATA_WIDTH-1:47*FORCE_DATA_WIDTH] = force_and_addr[46*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:46*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[48*FORCE_DATA_WIDTH-1:47*FORCE_DATA_WIDTH] = force_and_addr[47*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:47*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[48*FORCE_DATA_WIDTH-1:47*FORCE_DATA_WIDTH] = force_and_addr[48*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:48*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[48*FORCE_DATA_WIDTH-1:47*FORCE_DATA_WIDTH] = force_and_addr[56*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:56*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[48*FORCE_DATA_WIDTH-1:47*FORCE_DATA_WIDTH] = force_and_addr[59*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:59*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[48*FORCE_DATA_WIDTH-1:47*FORCE_DATA_WIDTH] = force_and_addr[60*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:60*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[48*FORCE_DATA_WIDTH-1:47*FORCE_DATA_WIDTH] = force_and_addr[62*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:62*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[48*FORCE_DATA_WIDTH-1:47*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[49*(NUM_NEIGHBOR_CELLS+1)-1:48*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[49*FORCE_DATA_WIDTH-1:48*FORCE_DATA_WIDTH] = force_and_addr[1*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:1*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[49*FORCE_DATA_WIDTH-1:48*FORCE_DATA_WIDTH] = force_and_addr[3*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:3*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[49*FORCE_DATA_WIDTH-1:48*FORCE_DATA_WIDTH] = force_and_addr[5*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:5*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[49*FORCE_DATA_WIDTH-1:48*FORCE_DATA_WIDTH] = force_and_addr[12*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:12*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[49*FORCE_DATA_WIDTH-1:48*FORCE_DATA_WIDTH] = force_and_addr[13*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:13*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[49*FORCE_DATA_WIDTH-1:48*FORCE_DATA_WIDTH] = force_and_addr[32*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:32*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[49*FORCE_DATA_WIDTH-1:48*FORCE_DATA_WIDTH] = force_and_addr[37*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:37*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[49*FORCE_DATA_WIDTH-1:48*FORCE_DATA_WIDTH] = force_and_addr[44*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:44*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[49*FORCE_DATA_WIDTH-1:48*FORCE_DATA_WIDTH] = force_and_addr[45*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:45*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[49*FORCE_DATA_WIDTH-1:48*FORCE_DATA_WIDTH] = force_and_addr[48*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:48*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[49*FORCE_DATA_WIDTH-1:48*FORCE_DATA_WIDTH] = force_and_addr[51*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:51*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[49*FORCE_DATA_WIDTH-1:48*FORCE_DATA_WIDTH] = force_and_addr[52*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:52*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[49*FORCE_DATA_WIDTH-1:48*FORCE_DATA_WIDTH] = force_and_addr[53*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:53*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[49*FORCE_DATA_WIDTH-1:48*FORCE_DATA_WIDTH] = force_and_addr[61*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:61*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[49*FORCE_DATA_WIDTH-1:48*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[50*(NUM_NEIGHBOR_CELLS+1)-1:49*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[50*FORCE_DATA_WIDTH-1:49*FORCE_DATA_WIDTH] = force_and_addr[0*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:0*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[50*FORCE_DATA_WIDTH-1:49*FORCE_DATA_WIDTH] = force_and_addr[2*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:2*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[50*FORCE_DATA_WIDTH-1:49*FORCE_DATA_WIDTH] = force_and_addr[6*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:6*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[50*FORCE_DATA_WIDTH-1:49*FORCE_DATA_WIDTH] = force_and_addr[13*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:13*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[50*FORCE_DATA_WIDTH-1:49*FORCE_DATA_WIDTH] = force_and_addr[14*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:14*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[50*FORCE_DATA_WIDTH-1:49*FORCE_DATA_WIDTH] = force_and_addr[33*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:33*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[50*FORCE_DATA_WIDTH-1:49*FORCE_DATA_WIDTH] = force_and_addr[38*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:38*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[50*FORCE_DATA_WIDTH-1:49*FORCE_DATA_WIDTH] = force_and_addr[45*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:45*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[50*FORCE_DATA_WIDTH-1:49*FORCE_DATA_WIDTH] = force_and_addr[46*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:46*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[50*FORCE_DATA_WIDTH-1:49*FORCE_DATA_WIDTH] = force_and_addr[48*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:48*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[50*FORCE_DATA_WIDTH-1:49*FORCE_DATA_WIDTH] = force_and_addr[49*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:49*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[50*FORCE_DATA_WIDTH-1:49*FORCE_DATA_WIDTH] = force_and_addr[53*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:53*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[50*FORCE_DATA_WIDTH-1:49*FORCE_DATA_WIDTH] = force_and_addr[54*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:54*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[50*FORCE_DATA_WIDTH-1:49*FORCE_DATA_WIDTH] = force_and_addr[62*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:62*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[50*FORCE_DATA_WIDTH-1:49*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[51*(NUM_NEIGHBOR_CELLS+1)-1:50*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[51*FORCE_DATA_WIDTH-1:50*FORCE_DATA_WIDTH] = force_and_addr[1*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:1*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[51*FORCE_DATA_WIDTH-1:50*FORCE_DATA_WIDTH] = force_and_addr[3*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:3*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[51*FORCE_DATA_WIDTH-1:50*FORCE_DATA_WIDTH] = force_and_addr[7*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:7*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[51*FORCE_DATA_WIDTH-1:50*FORCE_DATA_WIDTH] = force_and_addr[14*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:14*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[51*FORCE_DATA_WIDTH-1:50*FORCE_DATA_WIDTH] = force_and_addr[15*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:15*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[51*FORCE_DATA_WIDTH-1:50*FORCE_DATA_WIDTH] = force_and_addr[34*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:34*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[51*FORCE_DATA_WIDTH-1:50*FORCE_DATA_WIDTH] = force_and_addr[39*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:39*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[51*FORCE_DATA_WIDTH-1:50*FORCE_DATA_WIDTH] = force_and_addr[46*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:46*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[51*FORCE_DATA_WIDTH-1:50*FORCE_DATA_WIDTH] = force_and_addr[47*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:47*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[51*FORCE_DATA_WIDTH-1:50*FORCE_DATA_WIDTH] = force_and_addr[49*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:49*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[51*FORCE_DATA_WIDTH-1:50*FORCE_DATA_WIDTH] = force_and_addr[50*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:50*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[51*FORCE_DATA_WIDTH-1:50*FORCE_DATA_WIDTH] = force_and_addr[54*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:54*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[51*FORCE_DATA_WIDTH-1:50*FORCE_DATA_WIDTH] = force_and_addr[55*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:55*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[51*FORCE_DATA_WIDTH-1:50*FORCE_DATA_WIDTH] = force_and_addr[63*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:63*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[51*FORCE_DATA_WIDTH-1:50*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[52*(NUM_NEIGHBOR_CELLS+1)-1:51*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[52*FORCE_DATA_WIDTH-1:51*FORCE_DATA_WIDTH] = force_and_addr[0*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:0*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[52*FORCE_DATA_WIDTH-1:51*FORCE_DATA_WIDTH] = force_and_addr[2*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:2*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[52*FORCE_DATA_WIDTH-1:51*FORCE_DATA_WIDTH] = force_and_addr[4*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:4*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[52*FORCE_DATA_WIDTH-1:51*FORCE_DATA_WIDTH] = force_and_addr[12*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:12*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[52*FORCE_DATA_WIDTH-1:51*FORCE_DATA_WIDTH] = force_and_addr[15*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:15*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[52*FORCE_DATA_WIDTH-1:51*FORCE_DATA_WIDTH] = force_and_addr[35*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:35*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[52*FORCE_DATA_WIDTH-1:51*FORCE_DATA_WIDTH] = force_and_addr[36*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:36*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[52*FORCE_DATA_WIDTH-1:51*FORCE_DATA_WIDTH] = force_and_addr[44*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:44*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[52*FORCE_DATA_WIDTH-1:51*FORCE_DATA_WIDTH] = force_and_addr[47*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:47*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[52*FORCE_DATA_WIDTH-1:51*FORCE_DATA_WIDTH] = force_and_addr[50*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:50*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[52*FORCE_DATA_WIDTH-1:51*FORCE_DATA_WIDTH] = force_and_addr[51*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:51*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[52*FORCE_DATA_WIDTH-1:51*FORCE_DATA_WIDTH] = force_and_addr[52*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:52*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[52*FORCE_DATA_WIDTH-1:51*FORCE_DATA_WIDTH] = force_and_addr[55*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:55*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[52*FORCE_DATA_WIDTH-1:51*FORCE_DATA_WIDTH] = force_and_addr[60*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:60*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[52*FORCE_DATA_WIDTH-1:51*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[53*(NUM_NEIGHBOR_CELLS+1)-1:52*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[53*FORCE_DATA_WIDTH-1:52*FORCE_DATA_WIDTH] = force_and_addr[0*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:0*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[53*FORCE_DATA_WIDTH-1:52*FORCE_DATA_WIDTH] = force_and_addr[1*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:1*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[53*FORCE_DATA_WIDTH-1:52*FORCE_DATA_WIDTH] = force_and_addr[5*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:5*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[53*FORCE_DATA_WIDTH-1:52*FORCE_DATA_WIDTH] = force_and_addr[7*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:7*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[53*FORCE_DATA_WIDTH-1:52*FORCE_DATA_WIDTH] = force_and_addr[9*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:9*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[53*FORCE_DATA_WIDTH-1:52*FORCE_DATA_WIDTH] = force_and_addr[32*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:32*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[53*FORCE_DATA_WIDTH-1:52*FORCE_DATA_WIDTH] = force_and_addr[33*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:33*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[53*FORCE_DATA_WIDTH-1:52*FORCE_DATA_WIDTH] = force_and_addr[36*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:36*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[53*FORCE_DATA_WIDTH-1:52*FORCE_DATA_WIDTH] = force_and_addr[41*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:41*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[53*FORCE_DATA_WIDTH-1:52*FORCE_DATA_WIDTH] = force_and_addr[49*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:49*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[53*FORCE_DATA_WIDTH-1:52*FORCE_DATA_WIDTH] = force_and_addr[52*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:52*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[53*FORCE_DATA_WIDTH-1:52*FORCE_DATA_WIDTH] = force_and_addr[55*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:55*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[53*FORCE_DATA_WIDTH-1:52*FORCE_DATA_WIDTH] = force_and_addr[56*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:56*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[53*FORCE_DATA_WIDTH-1:52*FORCE_DATA_WIDTH] = force_and_addr[57*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:57*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[53*FORCE_DATA_WIDTH-1:52*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[54*(NUM_NEIGHBOR_CELLS+1)-1:53*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[54*FORCE_DATA_WIDTH-1:53*FORCE_DATA_WIDTH] = force_and_addr[1*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:1*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[54*FORCE_DATA_WIDTH-1:53*FORCE_DATA_WIDTH] = force_and_addr[2*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:2*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[54*FORCE_DATA_WIDTH-1:53*FORCE_DATA_WIDTH] = force_and_addr[4*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:4*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[54*FORCE_DATA_WIDTH-1:53*FORCE_DATA_WIDTH] = force_and_addr[6*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:6*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[54*FORCE_DATA_WIDTH-1:53*FORCE_DATA_WIDTH] = force_and_addr[10*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:10*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[54*FORCE_DATA_WIDTH-1:53*FORCE_DATA_WIDTH] = force_and_addr[33*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:33*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[54*FORCE_DATA_WIDTH-1:53*FORCE_DATA_WIDTH] = force_and_addr[34*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:34*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[54*FORCE_DATA_WIDTH-1:53*FORCE_DATA_WIDTH] = force_and_addr[37*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:37*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[54*FORCE_DATA_WIDTH-1:53*FORCE_DATA_WIDTH] = force_and_addr[42*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:42*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[54*FORCE_DATA_WIDTH-1:53*FORCE_DATA_WIDTH] = force_and_addr[50*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:50*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[54*FORCE_DATA_WIDTH-1:53*FORCE_DATA_WIDTH] = force_and_addr[52*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:52*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[54*FORCE_DATA_WIDTH-1:53*FORCE_DATA_WIDTH] = force_and_addr[53*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:53*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[54*FORCE_DATA_WIDTH-1:53*FORCE_DATA_WIDTH] = force_and_addr[57*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:57*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[54*FORCE_DATA_WIDTH-1:53*FORCE_DATA_WIDTH] = force_and_addr[58*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:58*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[54*FORCE_DATA_WIDTH-1:53*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[55*(NUM_NEIGHBOR_CELLS+1)-1:54*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[55*FORCE_DATA_WIDTH-1:54*FORCE_DATA_WIDTH] = force_and_addr[2*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:2*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[55*FORCE_DATA_WIDTH-1:54*FORCE_DATA_WIDTH] = force_and_addr[3*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:3*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[55*FORCE_DATA_WIDTH-1:54*FORCE_DATA_WIDTH] = force_and_addr[5*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:5*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[55*FORCE_DATA_WIDTH-1:54*FORCE_DATA_WIDTH] = force_and_addr[7*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:7*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[55*FORCE_DATA_WIDTH-1:54*FORCE_DATA_WIDTH] = force_and_addr[11*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:11*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[55*FORCE_DATA_WIDTH-1:54*FORCE_DATA_WIDTH] = force_and_addr[34*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:34*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[55*FORCE_DATA_WIDTH-1:54*FORCE_DATA_WIDTH] = force_and_addr[35*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:35*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[55*FORCE_DATA_WIDTH-1:54*FORCE_DATA_WIDTH] = force_and_addr[38*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:38*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[55*FORCE_DATA_WIDTH-1:54*FORCE_DATA_WIDTH] = force_and_addr[43*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:43*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[55*FORCE_DATA_WIDTH-1:54*FORCE_DATA_WIDTH] = force_and_addr[51*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:51*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[55*FORCE_DATA_WIDTH-1:54*FORCE_DATA_WIDTH] = force_and_addr[53*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:53*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[55*FORCE_DATA_WIDTH-1:54*FORCE_DATA_WIDTH] = force_and_addr[54*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:54*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[55*FORCE_DATA_WIDTH-1:54*FORCE_DATA_WIDTH] = force_and_addr[58*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:58*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[55*FORCE_DATA_WIDTH-1:54*FORCE_DATA_WIDTH] = force_and_addr[59*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:59*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[55*FORCE_DATA_WIDTH-1:54*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[56*(NUM_NEIGHBOR_CELLS+1)-1:55*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[56*FORCE_DATA_WIDTH-1:55*FORCE_DATA_WIDTH] = force_and_addr[0*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:0*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[56*FORCE_DATA_WIDTH-1:55*FORCE_DATA_WIDTH] = force_and_addr[3*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:3*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[56*FORCE_DATA_WIDTH-1:55*FORCE_DATA_WIDTH] = force_and_addr[4*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:4*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[56*FORCE_DATA_WIDTH-1:55*FORCE_DATA_WIDTH] = force_and_addr[6*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:6*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[56*FORCE_DATA_WIDTH-1:55*FORCE_DATA_WIDTH] = force_and_addr[8*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:8*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[56*FORCE_DATA_WIDTH-1:55*FORCE_DATA_WIDTH] = force_and_addr[32*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:32*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[56*FORCE_DATA_WIDTH-1:55*FORCE_DATA_WIDTH] = force_and_addr[35*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:35*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[56*FORCE_DATA_WIDTH-1:55*FORCE_DATA_WIDTH] = force_and_addr[39*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:39*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[56*FORCE_DATA_WIDTH-1:55*FORCE_DATA_WIDTH] = force_and_addr[40*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:40*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[56*FORCE_DATA_WIDTH-1:55*FORCE_DATA_WIDTH] = force_and_addr[48*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:48*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[56*FORCE_DATA_WIDTH-1:55*FORCE_DATA_WIDTH] = force_and_addr[54*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:54*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[56*FORCE_DATA_WIDTH-1:55*FORCE_DATA_WIDTH] = force_and_addr[55*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:55*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[56*FORCE_DATA_WIDTH-1:55*FORCE_DATA_WIDTH] = force_and_addr[56*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:56*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[56*FORCE_DATA_WIDTH-1:55*FORCE_DATA_WIDTH] = force_and_addr[59*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:59*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[56*FORCE_DATA_WIDTH-1:55*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[57*(NUM_NEIGHBOR_CELLS+1)-1:56*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[57*FORCE_DATA_WIDTH-1:56*FORCE_DATA_WIDTH] = force_and_addr[4*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:4*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[57*FORCE_DATA_WIDTH-1:56*FORCE_DATA_WIDTH] = force_and_addr[5*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:5*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[57*FORCE_DATA_WIDTH-1:56*FORCE_DATA_WIDTH] = force_and_addr[9*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:9*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[57*FORCE_DATA_WIDTH-1:56*FORCE_DATA_WIDTH] = force_and_addr[11*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:11*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[57*FORCE_DATA_WIDTH-1:56*FORCE_DATA_WIDTH] = force_and_addr[13*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:13*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[57*FORCE_DATA_WIDTH-1:56*FORCE_DATA_WIDTH] = force_and_addr[36*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:36*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[57*FORCE_DATA_WIDTH-1:56*FORCE_DATA_WIDTH] = force_and_addr[37*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:37*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[57*FORCE_DATA_WIDTH-1:56*FORCE_DATA_WIDTH] = force_and_addr[40*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:40*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[57*FORCE_DATA_WIDTH-1:56*FORCE_DATA_WIDTH] = force_and_addr[45*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:45*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[57*FORCE_DATA_WIDTH-1:56*FORCE_DATA_WIDTH] = force_and_addr[53*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:53*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[57*FORCE_DATA_WIDTH-1:56*FORCE_DATA_WIDTH] = force_and_addr[56*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:56*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[57*FORCE_DATA_WIDTH-1:56*FORCE_DATA_WIDTH] = force_and_addr[59*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:59*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[57*FORCE_DATA_WIDTH-1:56*FORCE_DATA_WIDTH] = force_and_addr[60*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:60*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[57*FORCE_DATA_WIDTH-1:56*FORCE_DATA_WIDTH] = force_and_addr[61*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:61*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[57*FORCE_DATA_WIDTH-1:56*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[58*(NUM_NEIGHBOR_CELLS+1)-1:57*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[58*FORCE_DATA_WIDTH-1:57*FORCE_DATA_WIDTH] = force_and_addr[5*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:5*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[58*FORCE_DATA_WIDTH-1:57*FORCE_DATA_WIDTH] = force_and_addr[6*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:6*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[58*FORCE_DATA_WIDTH-1:57*FORCE_DATA_WIDTH] = force_and_addr[8*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:8*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[58*FORCE_DATA_WIDTH-1:57*FORCE_DATA_WIDTH] = force_and_addr[10*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:10*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[58*FORCE_DATA_WIDTH-1:57*FORCE_DATA_WIDTH] = force_and_addr[14*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:14*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[58*FORCE_DATA_WIDTH-1:57*FORCE_DATA_WIDTH] = force_and_addr[37*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:37*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[58*FORCE_DATA_WIDTH-1:57*FORCE_DATA_WIDTH] = force_and_addr[38*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:38*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[58*FORCE_DATA_WIDTH-1:57*FORCE_DATA_WIDTH] = force_and_addr[41*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:41*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[58*FORCE_DATA_WIDTH-1:57*FORCE_DATA_WIDTH] = force_and_addr[46*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:46*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[58*FORCE_DATA_WIDTH-1:57*FORCE_DATA_WIDTH] = force_and_addr[54*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:54*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[58*FORCE_DATA_WIDTH-1:57*FORCE_DATA_WIDTH] = force_and_addr[56*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:56*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[58*FORCE_DATA_WIDTH-1:57*FORCE_DATA_WIDTH] = force_and_addr[57*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:57*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[58*FORCE_DATA_WIDTH-1:57*FORCE_DATA_WIDTH] = force_and_addr[61*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:61*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[58*FORCE_DATA_WIDTH-1:57*FORCE_DATA_WIDTH] = force_and_addr[62*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:62*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[58*FORCE_DATA_WIDTH-1:57*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[59*(NUM_NEIGHBOR_CELLS+1)-1:58*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[59*FORCE_DATA_WIDTH-1:58*FORCE_DATA_WIDTH] = force_and_addr[6*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:6*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[59*FORCE_DATA_WIDTH-1:58*FORCE_DATA_WIDTH] = force_and_addr[7*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:7*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[59*FORCE_DATA_WIDTH-1:58*FORCE_DATA_WIDTH] = force_and_addr[9*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:9*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[59*FORCE_DATA_WIDTH-1:58*FORCE_DATA_WIDTH] = force_and_addr[11*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:11*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[59*FORCE_DATA_WIDTH-1:58*FORCE_DATA_WIDTH] = force_and_addr[15*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:15*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[59*FORCE_DATA_WIDTH-1:58*FORCE_DATA_WIDTH] = force_and_addr[38*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:38*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[59*FORCE_DATA_WIDTH-1:58*FORCE_DATA_WIDTH] = force_and_addr[39*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:39*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[59*FORCE_DATA_WIDTH-1:58*FORCE_DATA_WIDTH] = force_and_addr[42*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:42*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[59*FORCE_DATA_WIDTH-1:58*FORCE_DATA_WIDTH] = force_and_addr[47*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:47*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[59*FORCE_DATA_WIDTH-1:58*FORCE_DATA_WIDTH] = force_and_addr[55*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:55*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[59*FORCE_DATA_WIDTH-1:58*FORCE_DATA_WIDTH] = force_and_addr[57*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:57*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[59*FORCE_DATA_WIDTH-1:58*FORCE_DATA_WIDTH] = force_and_addr[58*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:58*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[59*FORCE_DATA_WIDTH-1:58*FORCE_DATA_WIDTH] = force_and_addr[62*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:62*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[59*FORCE_DATA_WIDTH-1:58*FORCE_DATA_WIDTH] = force_and_addr[63*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:63*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[59*FORCE_DATA_WIDTH-1:58*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[60*(NUM_NEIGHBOR_CELLS+1)-1:59*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[60*FORCE_DATA_WIDTH-1:59*FORCE_DATA_WIDTH] = force_and_addr[4*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:4*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[60*FORCE_DATA_WIDTH-1:59*FORCE_DATA_WIDTH] = force_and_addr[7*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:7*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[60*FORCE_DATA_WIDTH-1:59*FORCE_DATA_WIDTH] = force_and_addr[8*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:8*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[60*FORCE_DATA_WIDTH-1:59*FORCE_DATA_WIDTH] = force_and_addr[10*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:10*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[60*FORCE_DATA_WIDTH-1:59*FORCE_DATA_WIDTH] = force_and_addr[12*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:12*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[60*FORCE_DATA_WIDTH-1:59*FORCE_DATA_WIDTH] = force_and_addr[36*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:36*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[60*FORCE_DATA_WIDTH-1:59*FORCE_DATA_WIDTH] = force_and_addr[39*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:39*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[60*FORCE_DATA_WIDTH-1:59*FORCE_DATA_WIDTH] = force_and_addr[43*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:43*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[60*FORCE_DATA_WIDTH-1:59*FORCE_DATA_WIDTH] = force_and_addr[44*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:44*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[60*FORCE_DATA_WIDTH-1:59*FORCE_DATA_WIDTH] = force_and_addr[52*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:52*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[60*FORCE_DATA_WIDTH-1:59*FORCE_DATA_WIDTH] = force_and_addr[58*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:58*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[60*FORCE_DATA_WIDTH-1:59*FORCE_DATA_WIDTH] = force_and_addr[59*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:59*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[60*FORCE_DATA_WIDTH-1:59*FORCE_DATA_WIDTH] = force_and_addr[60*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:60*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[60*FORCE_DATA_WIDTH-1:59*FORCE_DATA_WIDTH] = force_and_addr[63*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:63*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[60*FORCE_DATA_WIDTH-1:59*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[61*(NUM_NEIGHBOR_CELLS+1)-1:60*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[61*FORCE_DATA_WIDTH-1:60*FORCE_DATA_WIDTH] = force_and_addr[1*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:1*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[61*FORCE_DATA_WIDTH-1:60*FORCE_DATA_WIDTH] = force_and_addr[8*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:8*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[61*FORCE_DATA_WIDTH-1:60*FORCE_DATA_WIDTH] = force_and_addr[9*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:9*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[61*FORCE_DATA_WIDTH-1:60*FORCE_DATA_WIDTH] = force_and_addr[13*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:13*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[61*FORCE_DATA_WIDTH-1:60*FORCE_DATA_WIDTH] = force_and_addr[15*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:15*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[61*FORCE_DATA_WIDTH-1:60*FORCE_DATA_WIDTH] = force_and_addr[33*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:33*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[61*FORCE_DATA_WIDTH-1:60*FORCE_DATA_WIDTH] = force_and_addr[40*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:40*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[61*FORCE_DATA_WIDTH-1:60*FORCE_DATA_WIDTH] = force_and_addr[41*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:41*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[61*FORCE_DATA_WIDTH-1:60*FORCE_DATA_WIDTH] = force_and_addr[44*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:44*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[61*FORCE_DATA_WIDTH-1:60*FORCE_DATA_WIDTH] = force_and_addr[48*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:48*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[61*FORCE_DATA_WIDTH-1:60*FORCE_DATA_WIDTH] = force_and_addr[49*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:49*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[61*FORCE_DATA_WIDTH-1:60*FORCE_DATA_WIDTH] = force_and_addr[57*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:57*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[61*FORCE_DATA_WIDTH-1:60*FORCE_DATA_WIDTH] = force_and_addr[60*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:60*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[61*FORCE_DATA_WIDTH-1:60*FORCE_DATA_WIDTH] = force_and_addr[63*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:63*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[61*FORCE_DATA_WIDTH-1:60*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[62*(NUM_NEIGHBOR_CELLS+1)-1:61*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[62*FORCE_DATA_WIDTH-1:61*FORCE_DATA_WIDTH] = force_and_addr[2*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:2*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[62*FORCE_DATA_WIDTH-1:61*FORCE_DATA_WIDTH] = force_and_addr[9*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:9*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[62*FORCE_DATA_WIDTH-1:61*FORCE_DATA_WIDTH] = force_and_addr[10*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:10*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[62*FORCE_DATA_WIDTH-1:61*FORCE_DATA_WIDTH] = force_and_addr[12*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:12*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[62*FORCE_DATA_WIDTH-1:61*FORCE_DATA_WIDTH] = force_and_addr[14*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:14*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[62*FORCE_DATA_WIDTH-1:61*FORCE_DATA_WIDTH] = force_and_addr[34*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:34*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[62*FORCE_DATA_WIDTH-1:61*FORCE_DATA_WIDTH] = force_and_addr[41*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:41*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[62*FORCE_DATA_WIDTH-1:61*FORCE_DATA_WIDTH] = force_and_addr[42*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:42*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[62*FORCE_DATA_WIDTH-1:61*FORCE_DATA_WIDTH] = force_and_addr[45*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:45*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[62*FORCE_DATA_WIDTH-1:61*FORCE_DATA_WIDTH] = force_and_addr[49*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:49*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[62*FORCE_DATA_WIDTH-1:61*FORCE_DATA_WIDTH] = force_and_addr[50*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:50*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[62*FORCE_DATA_WIDTH-1:61*FORCE_DATA_WIDTH] = force_and_addr[58*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:58*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[62*FORCE_DATA_WIDTH-1:61*FORCE_DATA_WIDTH] = force_and_addr[60*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:60*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[62*FORCE_DATA_WIDTH-1:61*FORCE_DATA_WIDTH] = force_and_addr[61*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:61*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[62*FORCE_DATA_WIDTH-1:61*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[63*(NUM_NEIGHBOR_CELLS+1)-1:62*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[63*FORCE_DATA_WIDTH-1:62*FORCE_DATA_WIDTH] = force_and_addr[3*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:3*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[63*FORCE_DATA_WIDTH-1:62*FORCE_DATA_WIDTH] = force_and_addr[10*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:10*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[63*FORCE_DATA_WIDTH-1:62*FORCE_DATA_WIDTH] = force_and_addr[11*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:11*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[63*FORCE_DATA_WIDTH-1:62*FORCE_DATA_WIDTH] = force_and_addr[13*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:13*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[63*FORCE_DATA_WIDTH-1:62*FORCE_DATA_WIDTH] = force_and_addr[15*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:15*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[63*FORCE_DATA_WIDTH-1:62*FORCE_DATA_WIDTH] = force_and_addr[35*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:35*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[63*FORCE_DATA_WIDTH-1:62*FORCE_DATA_WIDTH] = force_and_addr[42*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:42*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[63*FORCE_DATA_WIDTH-1:62*FORCE_DATA_WIDTH] = force_and_addr[43*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:43*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[63*FORCE_DATA_WIDTH-1:62*FORCE_DATA_WIDTH] = force_and_addr[46*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:46*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[63*FORCE_DATA_WIDTH-1:62*FORCE_DATA_WIDTH] = force_and_addr[50*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:50*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[63*FORCE_DATA_WIDTH-1:62*FORCE_DATA_WIDTH] = force_and_addr[51*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:51*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[63*FORCE_DATA_WIDTH-1:62*FORCE_DATA_WIDTH] = force_and_addr[59*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:59*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[63*FORCE_DATA_WIDTH-1:62*FORCE_DATA_WIDTH] = force_and_addr[61*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:61*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[63*FORCE_DATA_WIDTH-1:62*FORCE_DATA_WIDTH] = force_and_addr[62*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:62*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[63*FORCE_DATA_WIDTH-1:62*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end
always@(*)
	begin
	case(arbitration_result[64*(NUM_NEIGHBOR_CELLS+1)-1:63*(NUM_NEIGHBOR_CELLS+1)])
		14'b00000000000001: 
			begin
			force_to_caches[64*FORCE_DATA_WIDTH-1:63*FORCE_DATA_WIDTH] = force_and_addr[0*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:0*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		14'b00000000000010: 
			begin
			force_to_caches[64*FORCE_DATA_WIDTH-1:63*FORCE_DATA_WIDTH] = force_and_addr[8*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:8*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00000000000100: 
			begin
			force_to_caches[64*FORCE_DATA_WIDTH-1:63*FORCE_DATA_WIDTH] = force_and_addr[11*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:11*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00000000001000: 
			begin
			force_to_caches[64*FORCE_DATA_WIDTH-1:63*FORCE_DATA_WIDTH] = force_and_addr[12*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:12*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000010000: 
			begin
			force_to_caches[64*FORCE_DATA_WIDTH-1:63*FORCE_DATA_WIDTH] = force_and_addr[14*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH-1:14*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH];
			end
		14'b00000000100000: 
			begin
			force_to_caches[64*FORCE_DATA_WIDTH-1:63*FORCE_DATA_WIDTH] = force_and_addr[32*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:32*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b00000001000000: 
			begin
			force_to_caches[64*FORCE_DATA_WIDTH-1:63*FORCE_DATA_WIDTH] = force_and_addr[40*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:40*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00000010000000: 
			begin
			force_to_caches[64*FORCE_DATA_WIDTH-1:63*FORCE_DATA_WIDTH] = force_and_addr[43*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:43*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b00000100000000: 
			begin
			force_to_caches[64*FORCE_DATA_WIDTH-1:63*FORCE_DATA_WIDTH] = force_and_addr[47*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH-1:47*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH];
			end
		14'b00001000000000: 
			begin
			force_to_caches[64*FORCE_DATA_WIDTH-1:63*FORCE_DATA_WIDTH] = force_and_addr[48*NUM_FILTER*FORCE_DATA_WIDTH+4*FORCE_DATA_WIDTH-1:48*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH];
			end
		14'b00010000000000: 
			begin
			force_to_caches[64*FORCE_DATA_WIDTH-1:63*FORCE_DATA_WIDTH] = force_and_addr[51*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH-1:51*NUM_FILTER*FORCE_DATA_WIDTH+5*FORCE_DATA_WIDTH];
			end
		14'b00100000000000: 
			begin
			force_to_caches[64*FORCE_DATA_WIDTH-1:63*FORCE_DATA_WIDTH] = force_and_addr[56*NUM_FILTER*FORCE_DATA_WIDTH+3*FORCE_DATA_WIDTH-1:56*NUM_FILTER*FORCE_DATA_WIDTH+2*FORCE_DATA_WIDTH];
			end
		14'b01000000000000: 
			begin
			force_to_caches[64*FORCE_DATA_WIDTH-1:63*FORCE_DATA_WIDTH] = force_and_addr[62*NUM_FILTER*FORCE_DATA_WIDTH+7*FORCE_DATA_WIDTH-1:62*NUM_FILTER*FORCE_DATA_WIDTH+6*FORCE_DATA_WIDTH];
			end
		14'b10000000000000: 
			begin
			force_to_caches[64*FORCE_DATA_WIDTH-1:63*FORCE_DATA_WIDTH] = force_and_addr[63*NUM_FILTER*FORCE_DATA_WIDTH+1*FORCE_DATA_WIDTH-1:63*NUM_FILTER*FORCE_DATA_WIDTH+0*FORCE_DATA_WIDTH];
			end
		default:
			begin
			force_to_caches[64*FORCE_DATA_WIDTH-1:63*FORCE_DATA_WIDTH] = 0;
			end
	endcase
	end

endmodule