// FP_ACC_Test.v

// Generated using ACDS version 18.0 219

`timescale 1 ps / 1 ps
module FP_ACC_Test (
		input  wire [31:0] ax,     //     ax.ax
		input  wire [31:0] ay,     //     ay.ay
		input  wire        clk,    //    clk.clk
		input  wire        clr,    //    clr.clr
		input  wire        ena,    //    ena.ena
		output wire [31:0] result  // result.result
	);

	FP_ACC_Test_altera_s10fpdsp_block_180_n4zfgua s10fpdsp_block_0 (
		.clk    (clk),    //   input,   width = 1,    clk.clk
		.ena    (ena),    //   input,   width = 1,    ena.ena
		.clr    (clr),    //   input,   width = 1,    clr.clr
		.result (result), //  output,  width = 32, result.result
		.ax     (ax),     //   input,  width = 32,     ax.ax
		.ay     (ay)      //   input,  width = 32,     ay.ay
	);

endmodule
