// eSRAM_test.v

// Generated using ACDS version 18.0 219

`timescale 1 ps / 1 ps
module eSRAM_test (
		input  wire [35:0] c0_data_0,       //  ram_input.s2c0_da_0
		input  wire [14:0] c0_rdaddress_0,  //           .s2c0_adrb_0
		input  wire        c0_rden_n_0,     //           .s2c0_meb_n_0
		input  wire        c0_sd_n_0,       //           .s2c0_sd_n_0
		input  wire [14:0] c0_wraddress_0,  //           .s2c0_adra_0
		input  wire        c0_wren_n_0,     //           .s2c0_mea_n_0
		input  wire [35:0] c1_data_0,       //           .s2c1_da_0
		input  wire [14:0] c1_rdaddress_0,  //           .s2c1_adrb_0
		input  wire        c1_rden_n_0,     //           .s2c1_meb_n_0
		input  wire        c1_sd_n_0,       //           .s2c1_sd_n_0
		input  wire [14:0] c1_wraddress_0,  //           .s2c1_adra_0
		input  wire        c1_wren_n_0,     //           .s2c1_mea_n_0
		input  wire [35:0] c2_data_0,       //           .s2c2_da_0
		input  wire [14:0] c2_rdaddress_0,  //           .s2c2_adrb_0
		input  wire        c2_rden_n_0,     //           .s2c2_meb_n_0
		input  wire        c2_sd_n_0,       //           .s2c2_sd_n_0
		input  wire [14:0] c2_wraddress_0,  //           .s2c2_adra_0
		input  wire        c2_wren_n_0,     //           .s2c2_mea_n_0
		input  wire        refclk,          //           .clock
		output wire [35:0] c0_q_0,          // ram_output.s2c0_qb_0
		output wire [35:0] c1_q_0,          //           .s2c1_qb_0
		output wire [35:0] c2_q_0,          //           .s2c2_qb_0
		output wire        esram2f_clk,     //           .esram2f_clk
		output wire        iopll_lock2core  //           .iopll_lock2core
	);

	eSRAM_test_esram_180_nuaykua #(
		.c0_address_width  (15),
		.c1_address_width  (15),
		.c2_address_width  (15),
		.c3_address_width  (11),
		.c4_address_width  (11),
		.c5_address_width  (11),
		.c6_address_width  (11),
		.c7_address_width  (11),
		.c0_data_width     (36),
		.c1_data_width     (36),
		.c2_data_width     (36),
		.c3_data_width     (72),
		.c4_data_width     (72),
		.c5_data_width     (72),
		.c6_data_width     (72),
		.c7_data_width     (72),
		.c0_disable        ("FALSE"),
		.c1_disable        ("FALSE"),
		.c2_disable        ("FALSE"),
		.c3_disable        ("TRUE"),
		.c4_disable        ("TRUE"),
		.c5_disable        ("TRUE"),
		.c6_disable        ("TRUE"),
		.c7_disable        ("TRUE"),
		.c0_bank_enable    ("C0_EN_10BANK"),
		.c1_bank_enable    ("C1_EN_10BANK"),
		.c2_bank_enable    ("C2_EN_10BANK"),
		.c3_bank_enable    ("C3_EN_0BANK"),
		.c4_bank_enable    ("C4_EN_0BANK"),
		.c5_bank_enable    ("C5_EN_0BANK"),
		.c6_bank_enable    ("C6_EN_0BANK"),
		.c7_bank_enable    ("C7_EN_0BANK"),
		.c0_ecc_enable     ("FALSE"),
		.c1_ecc_enable     ("FALSE"),
		.c2_ecc_enable     ("FALSE"),
		.c3_ecc_enable     ("FALSE"),
		.c4_ecc_enable     ("FALSE"),
		.c5_ecc_enable     ("FALSE"),
		.c6_ecc_enable     ("FALSE"),
		.c7_ecc_enable     ("FALSE"),
		.c0_ecc_byp_enable ("FALSE"),
		.c1_ecc_byp_enable ("FALSE"),
		.c2_ecc_byp_enable ("FALSE"),
		.c3_ecc_byp_enable ("FALSE"),
		.c4_ecc_byp_enable ("FALSE"),
		.c5_ecc_byp_enable ("FALSE"),
		.c6_ecc_byp_enable ("FALSE"),
		.c7_ecc_byp_enable ("FALSE"),
		.c0_wr_fwd_enable  ("FALSE"),
		.c1_wr_fwd_enable  ("FALSE"),
		.c2_wr_fwd_enable  ("FALSE"),
		.c3_wr_fwd_enable  ("FALSE"),
		.c4_wr_fwd_enable  ("FALSE"),
		.c5_wr_fwd_enable  ("FALSE"),
		.c6_wr_fwd_enable  ("FALSE"),
		.c7_wr_fwd_enable  ("FALSE"),
		.c0_lpmode_enable  ("FALSE"),
		.c1_lpmode_enable  ("FALSE"),
		.c2_lpmode_enable  ("FALSE"),
		.c3_lpmode_enable  ("FALSE"),
		.c4_lpmode_enable  ("FALSE"),
		.c5_lpmode_enable  ("FALSE"),
		.c6_lpmode_enable  ("FALSE"),
		.c7_lpmode_enable  ("FALSE"),
		.clock_rate        ("FULLRATE")
	) esram_0 (
		.c0_q_0          (c0_q_0),          //  output,  width = 36, ram_output.s2c0_qb_0
		.c1_q_0          (c1_q_0),          //  output,  width = 36,           .s2c1_qb_0
		.c2_q_0          (c2_q_0),          //  output,  width = 36,           .s2c2_qb_0
		.esram2f_clk     (esram2f_clk),     //  output,   width = 1,           .esram2f_clk
		.iopll_lock2core (iopll_lock2core), //  output,   width = 1,           .iopll_lock2core
		.c0_data_0       (c0_data_0),       //   input,  width = 36,  ram_input.s2c0_da_0
		.c0_rdaddress_0  (c0_rdaddress_0),  //   input,  width = 15,           .s2c0_adrb_0
		.c0_rden_n_0     (c0_rden_n_0),     //   input,   width = 1,           .s2c0_meb_n_0
		.c0_sd_n_0       (c0_sd_n_0),       //   input,   width = 1,           .s2c0_sd_n_0
		.c0_wraddress_0  (c0_wraddress_0),  //   input,  width = 15,           .s2c0_adra_0
		.c0_wren_n_0     (c0_wren_n_0),     //   input,   width = 1,           .s2c0_mea_n_0
		.c1_data_0       (c1_data_0),       //   input,  width = 36,           .s2c1_da_0
		.c1_rdaddress_0  (c1_rdaddress_0),  //   input,  width = 15,           .s2c1_adrb_0
		.c1_rden_n_0     (c1_rden_n_0),     //   input,   width = 1,           .s2c1_meb_n_0
		.c1_sd_n_0       (c1_sd_n_0),       //   input,   width = 1,           .s2c1_sd_n_0
		.c1_wraddress_0  (c1_wraddress_0),  //   input,  width = 15,           .s2c1_adra_0
		.c1_wren_n_0     (c1_wren_n_0),     //   input,   width = 1,           .s2c1_mea_n_0
		.c2_data_0       (c2_data_0),       //   input,  width = 36,           .s2c2_da_0
		.c2_rdaddress_0  (c2_rdaddress_0),  //   input,  width = 15,           .s2c2_adrb_0
		.c2_rden_n_0     (c2_rden_n_0),     //   input,   width = 1,           .s2c2_meb_n_0
		.c2_sd_n_0       (c2_sd_n_0),       //   input,   width = 1,           .s2c2_sd_n_0
		.c2_wraddress_0  (c2_wraddress_0),  //   input,  width = 15,           .s2c2_adra_0
		.c2_wren_n_0     (c2_wren_n_0),     //   input,   width = 1,           .s2c2_mea_n_0
		.refclk          (refclk)           //   input,   width = 1,           .clock
	);

endmodule
