module FIX_SQRT (
		input  wire        clk,     //     clk.clk
		input  wire [0:0]  en,      //      en.en
		input  wire [31:0] radical, // radical.radical
		output wire [31:0] result,  //  result.result
		input  wire        rst      //     rst.reset
	);
endmodule

