module FP_GreaterThan_or_Equal (
		input  wire [31:0] a,      //      a.a
		input  wire        areset, // areset.reset
		input  wire [31:0] b,      //      b.b
		input  wire        clk,    //    clk.clk
		output wire [0:0]  q       //      q.q
	);
endmodule

