module arbitration_to_success_mapping
#(
	parameter NUM_CELLS = 64, 
	parameter NUM_NEIGHBOR_CELLS = 13, 
	parameter NUM_FILTER = 7
)
(
	input [NUM_CELLS*(NUM_NEIGHBOR_CELLS+1)-1:0] arbitration_result, 
	
	output [NUM_CELLS*NUM_FILTER-1:0] force_cache_write_success
);
assign force_cache_write_success[0] = arbitration_result[0*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[63*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[1] = arbitration_result[49*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[51*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[2] = arbitration_result[20*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[7*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[3] = arbitration_result[15*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[52*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[4] = arbitration_result[55*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[16*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[5] = arbitration_result[23*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[12*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[6] = arbitration_result[31*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[1*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[7] = arbitration_result[1*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[60*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[8] = arbitration_result[50*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[48*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[9] = arbitration_result[21*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[4*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[10] = arbitration_result[12*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[53*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[11] = arbitration_result[52*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[17*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[12] = arbitration_result[20*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[13*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[13] = arbitration_result[28*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[2*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[14] = arbitration_result[2*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[61*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[15] = arbitration_result[51*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[49*(NUM_NEIGHBOR_CELLS+1)+1];
assign force_cache_write_success[16] = arbitration_result[22*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[5*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[17] = arbitration_result[13*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[54*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[18] = arbitration_result[53*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[18*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[19] = arbitration_result[21*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[14*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[20] = arbitration_result[29*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[3*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[21] = arbitration_result[3*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[62*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[22] = arbitration_result[48*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[50*(NUM_NEIGHBOR_CELLS+1)+1];
assign force_cache_write_success[23] = arbitration_result[23*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[6*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[24] = arbitration_result[14*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[55*(NUM_NEIGHBOR_CELLS+1)+1];
assign force_cache_write_success[25] = arbitration_result[54*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[19*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[26] = arbitration_result[22*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[15*(NUM_NEIGHBOR_CELLS+1)+1];
assign force_cache_write_success[27] = arbitration_result[30*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[0*(NUM_NEIGHBOR_CELLS+1)+1];
assign force_cache_write_success[28] = arbitration_result[4*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[51*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[29] = arbitration_result[53*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[55*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[30] = arbitration_result[24*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[11*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[31] = arbitration_result[3*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[56*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[32] = arbitration_result[59*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[20*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[33] = arbitration_result[27*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[0*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[34] = arbitration_result[19*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[5*(NUM_NEIGHBOR_CELLS+1)+1];
assign force_cache_write_success[35] = arbitration_result[5*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[48*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[36] = arbitration_result[54*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[52*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[37] = arbitration_result[25*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[8*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[38] = arbitration_result[0*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[57*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[39] = arbitration_result[56*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[21*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[40] = arbitration_result[24*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[1*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[41] = arbitration_result[16*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[6*(NUM_NEIGHBOR_CELLS+1)+1];
assign force_cache_write_success[42] = arbitration_result[6*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[49*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[43] = arbitration_result[55*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[53*(NUM_NEIGHBOR_CELLS+1)+3];
assign force_cache_write_success[44] = arbitration_result[26*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[9*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[45] = arbitration_result[1*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[58*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[46] = arbitration_result[57*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[22*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[47] = arbitration_result[25*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[2*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[48] = arbitration_result[17*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[7*(NUM_NEIGHBOR_CELLS+1)+1];
assign force_cache_write_success[49] = arbitration_result[7*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[50*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[50] = arbitration_result[52*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[54*(NUM_NEIGHBOR_CELLS+1)+3];
assign force_cache_write_success[51] = arbitration_result[27*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[10*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[52] = arbitration_result[2*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[59*(NUM_NEIGHBOR_CELLS+1)+1];
assign force_cache_write_success[53] = arbitration_result[58*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[23*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[54] = arbitration_result[26*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[3*(NUM_NEIGHBOR_CELLS+1)+3];
assign force_cache_write_success[55] = arbitration_result[18*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[4*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[56] = arbitration_result[8*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[55*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[57] = arbitration_result[57*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[59*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[58] = arbitration_result[28*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[15*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[59] = arbitration_result[7*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[60*(NUM_NEIGHBOR_CELLS+1)+1];
assign force_cache_write_success[60] = arbitration_result[63*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[24*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[61] = arbitration_result[31*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[4*(NUM_NEIGHBOR_CELLS+1)+3];
assign force_cache_write_success[62] = arbitration_result[23*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[9*(NUM_NEIGHBOR_CELLS+1)+1];
assign force_cache_write_success[63] = arbitration_result[9*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[52*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[64] = arbitration_result[58*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[56*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[65] = arbitration_result[29*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[12*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[66] = arbitration_result[4*(NUM_NEIGHBOR_CELLS+1)+4] | arbitration_result[61*(NUM_NEIGHBOR_CELLS+1)+1];
assign force_cache_write_success[67] = arbitration_result[60*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[25*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[68] = arbitration_result[28*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[5*(NUM_NEIGHBOR_CELLS+1)+3];
assign force_cache_write_success[69] = arbitration_result[20*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[10*(NUM_NEIGHBOR_CELLS+1)+1];
assign force_cache_write_success[70] = arbitration_result[10*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[53*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[71] = arbitration_result[59*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[57*(NUM_NEIGHBOR_CELLS+1)+3];
assign force_cache_write_success[72] = arbitration_result[30*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[13*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[73] = arbitration_result[5*(NUM_NEIGHBOR_CELLS+1)+4] | arbitration_result[62*(NUM_NEIGHBOR_CELLS+1)+1];
assign force_cache_write_success[74] = arbitration_result[61*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[26*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[75] = arbitration_result[29*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[6*(NUM_NEIGHBOR_CELLS+1)+3];
assign force_cache_write_success[76] = arbitration_result[21*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[11*(NUM_NEIGHBOR_CELLS+1)+1];
assign force_cache_write_success[77] = arbitration_result[11*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[54*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[78] = arbitration_result[56*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[58*(NUM_NEIGHBOR_CELLS+1)+3];
assign force_cache_write_success[79] = arbitration_result[31*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[14*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[80] = arbitration_result[6*(NUM_NEIGHBOR_CELLS+1)+4] | arbitration_result[63*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[81] = arbitration_result[62*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[27*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[82] = arbitration_result[30*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[7*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[83] = arbitration_result[22*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[8*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[84] = arbitration_result[12*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[59*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[85] = arbitration_result[61*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[63*(NUM_NEIGHBOR_CELLS+1)+3];
assign force_cache_write_success[86] = arbitration_result[16*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[3*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[87] = arbitration_result[11*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[48*(NUM_NEIGHBOR_CELLS+1)+3];
assign force_cache_write_success[88] = arbitration_result[51*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[28*(NUM_NEIGHBOR_CELLS+1)+3];
assign force_cache_write_success[89] = arbitration_result[19*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[8*(NUM_NEIGHBOR_CELLS+1)+3];
assign force_cache_write_success[90] = arbitration_result[27*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[13*(NUM_NEIGHBOR_CELLS+1)+3];
assign force_cache_write_success[91] = arbitration_result[13*(NUM_NEIGHBOR_CELLS+1)+4] | arbitration_result[56*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[92] = arbitration_result[62*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[60*(NUM_NEIGHBOR_CELLS+1)+3];
assign force_cache_write_success[93] = arbitration_result[17*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[0*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[94] = arbitration_result[8*(NUM_NEIGHBOR_CELLS+1)+4] | arbitration_result[49*(NUM_NEIGHBOR_CELLS+1)+3];
assign force_cache_write_success[95] = arbitration_result[48*(NUM_NEIGHBOR_CELLS+1)+4] | arbitration_result[29*(NUM_NEIGHBOR_CELLS+1)+3];
assign force_cache_write_success[96] = arbitration_result[16*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[9*(NUM_NEIGHBOR_CELLS+1)+3];
assign force_cache_write_success[97] = arbitration_result[24*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[14*(NUM_NEIGHBOR_CELLS+1)+3];
assign force_cache_write_success[98] = arbitration_result[14*(NUM_NEIGHBOR_CELLS+1)+4] | arbitration_result[57*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[99] = arbitration_result[63*(NUM_NEIGHBOR_CELLS+1)+4] | arbitration_result[61*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[100] = arbitration_result[18*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[1*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[101] = arbitration_result[9*(NUM_NEIGHBOR_CELLS+1)+4] | arbitration_result[50*(NUM_NEIGHBOR_CELLS+1)+3];
assign force_cache_write_success[102] = arbitration_result[49*(NUM_NEIGHBOR_CELLS+1)+4] | arbitration_result[30*(NUM_NEIGHBOR_CELLS+1)+3];
assign force_cache_write_success[103] = arbitration_result[17*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[10*(NUM_NEIGHBOR_CELLS+1)+3];
assign force_cache_write_success[104] = arbitration_result[25*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[15*(NUM_NEIGHBOR_CELLS+1)+3];
assign force_cache_write_success[105] = arbitration_result[15*(NUM_NEIGHBOR_CELLS+1)+4] | arbitration_result[58*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[106] = arbitration_result[60*(NUM_NEIGHBOR_CELLS+1)+4] | arbitration_result[62*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[107] = arbitration_result[19*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[2*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[108] = arbitration_result[10*(NUM_NEIGHBOR_CELLS+1)+4] | arbitration_result[51*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[109] = arbitration_result[50*(NUM_NEIGHBOR_CELLS+1)+4] | arbitration_result[31*(NUM_NEIGHBOR_CELLS+1)+3];
assign force_cache_write_success[110] = arbitration_result[18*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[11*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[111] = arbitration_result[26*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[12*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[112] = arbitration_result[16*(NUM_NEIGHBOR_CELLS+1)+4] | arbitration_result[15*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[113] = arbitration_result[1*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[3*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[114] = arbitration_result[36*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[23*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[115] = arbitration_result[31*(NUM_NEIGHBOR_CELLS+1)+4] | arbitration_result[4*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[116] = arbitration_result[7*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[32*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[117] = arbitration_result[39*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[28*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[118] = arbitration_result[47*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[17*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[119] = arbitration_result[17*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[12*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[120] = arbitration_result[2*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[0*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[121] = arbitration_result[37*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[20*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[122] = arbitration_result[28*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[5*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[123] = arbitration_result[4*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[33*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[124] = arbitration_result[36*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[29*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[125] = arbitration_result[44*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[18*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[126] = arbitration_result[18*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[13*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[127] = arbitration_result[3*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[1*(NUM_NEIGHBOR_CELLS+1)+6];
assign force_cache_write_success[128] = arbitration_result[38*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[21*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[129] = arbitration_result[29*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[6*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[130] = arbitration_result[5*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[34*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[131] = arbitration_result[37*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[30*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[132] = arbitration_result[45*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[19*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[133] = arbitration_result[19*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[14*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[134] = arbitration_result[0*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[2*(NUM_NEIGHBOR_CELLS+1)+6];
assign force_cache_write_success[135] = arbitration_result[39*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[22*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[136] = arbitration_result[30*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[7*(NUM_NEIGHBOR_CELLS+1)+6];
assign force_cache_write_success[137] = arbitration_result[6*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[35*(NUM_NEIGHBOR_CELLS+1)+0];
assign force_cache_write_success[138] = arbitration_result[38*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[31*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[139] = arbitration_result[46*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[16*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[140] = arbitration_result[20*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[3*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[141] = arbitration_result[5*(NUM_NEIGHBOR_CELLS+1)+7] | arbitration_result[7*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[142] = arbitration_result[40*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[27*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[143] = arbitration_result[19*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[8*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[144] = arbitration_result[11*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[36*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[145] = arbitration_result[43*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[16*(NUM_NEIGHBOR_CELLS+1)+6];
assign force_cache_write_success[146] = arbitration_result[35*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[21*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[147] = arbitration_result[21*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[0*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[148] = arbitration_result[6*(NUM_NEIGHBOR_CELLS+1)+7] | arbitration_result[4*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[149] = arbitration_result[41*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[24*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[150] = arbitration_result[16*(NUM_NEIGHBOR_CELLS+1)+7] | arbitration_result[9*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[151] = arbitration_result[8*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[37*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[152] = arbitration_result[40*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[17*(NUM_NEIGHBOR_CELLS+1)+6];
assign force_cache_write_success[153] = arbitration_result[32*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[22*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[154] = arbitration_result[22*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[1*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[155] = arbitration_result[7*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[5*(NUM_NEIGHBOR_CELLS+1)+8];
assign force_cache_write_success[156] = arbitration_result[42*(NUM_NEIGHBOR_CELLS+1)+0] | arbitration_result[25*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[157] = arbitration_result[17*(NUM_NEIGHBOR_CELLS+1)+7] | arbitration_result[10*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[158] = arbitration_result[9*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[38*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[159] = arbitration_result[41*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[18*(NUM_NEIGHBOR_CELLS+1)+6];
assign force_cache_write_success[160] = arbitration_result[33*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[23*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[161] = arbitration_result[23*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[2*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[162] = arbitration_result[4*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[6*(NUM_NEIGHBOR_CELLS+1)+8];
assign force_cache_write_success[163] = arbitration_result[43*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[26*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[164] = arbitration_result[18*(NUM_NEIGHBOR_CELLS+1)+7] | arbitration_result[11*(NUM_NEIGHBOR_CELLS+1)+6];
assign force_cache_write_success[165] = arbitration_result[10*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[39*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[166] = arbitration_result[42*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[19*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[167] = arbitration_result[34*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[20*(NUM_NEIGHBOR_CELLS+1)+6];
assign force_cache_write_success[168] = arbitration_result[24*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[7*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[169] = arbitration_result[9*(NUM_NEIGHBOR_CELLS+1)+7] | arbitration_result[11*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[170] = arbitration_result[44*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[31*(NUM_NEIGHBOR_CELLS+1)+6];
assign force_cache_write_success[171] = arbitration_result[23*(NUM_NEIGHBOR_CELLS+1)+7] | arbitration_result[12*(NUM_NEIGHBOR_CELLS+1)+6];
assign force_cache_write_success[172] = arbitration_result[15*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[40*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[173] = arbitration_result[47*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[20*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[174] = arbitration_result[39*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[25*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[175] = arbitration_result[25*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[4*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[176] = arbitration_result[10*(NUM_NEIGHBOR_CELLS+1)+7] | arbitration_result[8*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[177] = arbitration_result[45*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[28*(NUM_NEIGHBOR_CELLS+1)+6];
assign force_cache_write_success[178] = arbitration_result[20*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[13*(NUM_NEIGHBOR_CELLS+1)+6];
assign force_cache_write_success[179] = arbitration_result[12*(NUM_NEIGHBOR_CELLS+1)+7] | arbitration_result[41*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[180] = arbitration_result[44*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[21*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[181] = arbitration_result[36*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[26*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[182] = arbitration_result[26*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[5*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[183] = arbitration_result[11*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[9*(NUM_NEIGHBOR_CELLS+1)+8];
assign force_cache_write_success[184] = arbitration_result[46*(NUM_NEIGHBOR_CELLS+1)+1] | arbitration_result[29*(NUM_NEIGHBOR_CELLS+1)+6];
assign force_cache_write_success[185] = arbitration_result[21*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[14*(NUM_NEIGHBOR_CELLS+1)+6];
assign force_cache_write_success[186] = arbitration_result[13*(NUM_NEIGHBOR_CELLS+1)+7] | arbitration_result[42*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[187] = arbitration_result[45*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[22*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[188] = arbitration_result[37*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[27*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[189] = arbitration_result[27*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[6*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[190] = arbitration_result[8*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[10*(NUM_NEIGHBOR_CELLS+1)+8];
assign force_cache_write_success[191] = arbitration_result[47*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[30*(NUM_NEIGHBOR_CELLS+1)+6];
assign force_cache_write_success[192] = arbitration_result[22*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[15*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[193] = arbitration_result[14*(NUM_NEIGHBOR_CELLS+1)+7] | arbitration_result[43*(NUM_NEIGHBOR_CELLS+1)+2];
assign force_cache_write_success[194] = arbitration_result[46*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[23*(NUM_NEIGHBOR_CELLS+1)+8];
assign force_cache_write_success[195] = arbitration_result[38*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[24*(NUM_NEIGHBOR_CELLS+1)+6];
assign force_cache_write_success[196] = arbitration_result[28*(NUM_NEIGHBOR_CELLS+1)+7] | arbitration_result[11*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[197] = arbitration_result[13*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[15*(NUM_NEIGHBOR_CELLS+1)+8];
assign force_cache_write_success[198] = arbitration_result[32*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[19*(NUM_NEIGHBOR_CELLS+1)+8];
assign force_cache_write_success[199] = arbitration_result[27*(NUM_NEIGHBOR_CELLS+1)+7] | arbitration_result[0*(NUM_NEIGHBOR_CELLS+1)+8];
assign force_cache_write_success[200] = arbitration_result[3*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[44*(NUM_NEIGHBOR_CELLS+1)+3];
assign force_cache_write_success[201] = arbitration_result[35*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[24*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[202] = arbitration_result[43*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[29*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[203] = arbitration_result[29*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[8*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[204] = arbitration_result[14*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[12*(NUM_NEIGHBOR_CELLS+1)+8];
assign force_cache_write_success[205] = arbitration_result[33*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[16*(NUM_NEIGHBOR_CELLS+1)+8];
assign force_cache_write_success[206] = arbitration_result[24*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[1*(NUM_NEIGHBOR_CELLS+1)+8];
assign force_cache_write_success[207] = arbitration_result[0*(NUM_NEIGHBOR_CELLS+1)+9] | arbitration_result[45*(NUM_NEIGHBOR_CELLS+1)+3];
assign force_cache_write_success[208] = arbitration_result[32*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[25*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[209] = arbitration_result[40*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[30*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[210] = arbitration_result[30*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[9*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[211] = arbitration_result[15*(NUM_NEIGHBOR_CELLS+1)+9] | arbitration_result[13*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[212] = arbitration_result[34*(NUM_NEIGHBOR_CELLS+1)+2] | arbitration_result[17*(NUM_NEIGHBOR_CELLS+1)+8];
assign force_cache_write_success[213] = arbitration_result[25*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[2*(NUM_NEIGHBOR_CELLS+1)+8];
assign force_cache_write_success[214] = arbitration_result[1*(NUM_NEIGHBOR_CELLS+1)+9] | arbitration_result[46*(NUM_NEIGHBOR_CELLS+1)+3];
assign force_cache_write_success[215] = arbitration_result[33*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[26*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[216] = arbitration_result[41*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[31*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[217] = arbitration_result[31*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[10*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[218] = arbitration_result[12*(NUM_NEIGHBOR_CELLS+1)+9] | arbitration_result[14*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[219] = arbitration_result[35*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[18*(NUM_NEIGHBOR_CELLS+1)+8];
assign force_cache_write_success[220] = arbitration_result[26*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[3*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[221] = arbitration_result[2*(NUM_NEIGHBOR_CELLS+1)+9] | arbitration_result[47*(NUM_NEIGHBOR_CELLS+1)+3];
assign force_cache_write_success[222] = arbitration_result[34*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[27*(NUM_NEIGHBOR_CELLS+1)+8];
assign force_cache_write_success[223] = arbitration_result[42*(NUM_NEIGHBOR_CELLS+1)+3] | arbitration_result[28*(NUM_NEIGHBOR_CELLS+1)+8];
assign force_cache_write_success[224] = arbitration_result[32*(NUM_NEIGHBOR_CELLS+1)+4] | arbitration_result[31*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[225] = arbitration_result[17*(NUM_NEIGHBOR_CELLS+1)+9] | arbitration_result[19*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[226] = arbitration_result[52*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[39*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[227] = arbitration_result[47*(NUM_NEIGHBOR_CELLS+1)+4] | arbitration_result[20*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[228] = arbitration_result[23*(NUM_NEIGHBOR_CELLS+1)+9] | arbitration_result[48*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[229] = arbitration_result[55*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[44*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[230] = arbitration_result[63*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[33*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[231] = arbitration_result[33*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[28*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[232] = arbitration_result[18*(NUM_NEIGHBOR_CELLS+1)+9] | arbitration_result[16*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[233] = arbitration_result[53*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[36*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[234] = arbitration_result[44*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[21*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[235] = arbitration_result[20*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[49*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[236] = arbitration_result[52*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[45*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[237] = arbitration_result[60*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[34*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[238] = arbitration_result[34*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[29*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[239] = arbitration_result[19*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[17*(NUM_NEIGHBOR_CELLS+1)+10];
assign force_cache_write_success[240] = arbitration_result[54*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[37*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[241] = arbitration_result[45*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[22*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[242] = arbitration_result[21*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[50*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[243] = arbitration_result[53*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[46*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[244] = arbitration_result[61*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[35*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[245] = arbitration_result[35*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[30*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[246] = arbitration_result[16*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[18*(NUM_NEIGHBOR_CELLS+1)+10];
assign force_cache_write_success[247] = arbitration_result[55*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[38*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[248] = arbitration_result[46*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[23*(NUM_NEIGHBOR_CELLS+1)+10];
assign force_cache_write_success[249] = arbitration_result[22*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[51*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[250] = arbitration_result[54*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[47*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[251] = arbitration_result[62*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[32*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[252] = arbitration_result[36*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[19*(NUM_NEIGHBOR_CELLS+1)+11];
assign force_cache_write_success[253] = arbitration_result[21*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[23*(NUM_NEIGHBOR_CELLS+1)+11];
assign force_cache_write_success[254] = arbitration_result[56*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[43*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[255] = arbitration_result[35*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[24*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[256] = arbitration_result[27*(NUM_NEIGHBOR_CELLS+1)+9] | arbitration_result[52*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[257] = arbitration_result[59*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[32*(NUM_NEIGHBOR_CELLS+1)+6];
assign force_cache_write_success[258] = arbitration_result[51*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[37*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[259] = arbitration_result[37*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[16*(NUM_NEIGHBOR_CELLS+1)+11];
assign force_cache_write_success[260] = arbitration_result[22*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[20*(NUM_NEIGHBOR_CELLS+1)+11];
assign force_cache_write_success[261] = arbitration_result[57*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[40*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[262] = arbitration_result[32*(NUM_NEIGHBOR_CELLS+1)+7] | arbitration_result[25*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[263] = arbitration_result[24*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[53*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[264] = arbitration_result[56*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[33*(NUM_NEIGHBOR_CELLS+1)+6];
assign force_cache_write_success[265] = arbitration_result[48*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[38*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[266] = arbitration_result[38*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[17*(NUM_NEIGHBOR_CELLS+1)+11];
assign force_cache_write_success[267] = arbitration_result[23*(NUM_NEIGHBOR_CELLS+1)+12] | arbitration_result[21*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[268] = arbitration_result[58*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[41*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[269] = arbitration_result[33*(NUM_NEIGHBOR_CELLS+1)+7] | arbitration_result[26*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[270] = arbitration_result[25*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[54*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[271] = arbitration_result[57*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[34*(NUM_NEIGHBOR_CELLS+1)+6];
assign force_cache_write_success[272] = arbitration_result[49*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[39*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[273] = arbitration_result[39*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[18*(NUM_NEIGHBOR_CELLS+1)+11];
assign force_cache_write_success[274] = arbitration_result[20*(NUM_NEIGHBOR_CELLS+1)+12] | arbitration_result[22*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[275] = arbitration_result[59*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[42*(NUM_NEIGHBOR_CELLS+1)+4];
assign force_cache_write_success[276] = arbitration_result[34*(NUM_NEIGHBOR_CELLS+1)+7] | arbitration_result[27*(NUM_NEIGHBOR_CELLS+1)+10];
assign force_cache_write_success[277] = arbitration_result[26*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[55*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[278] = arbitration_result[58*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[35*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[279] = arbitration_result[50*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[36*(NUM_NEIGHBOR_CELLS+1)+6];
assign force_cache_write_success[280] = arbitration_result[40*(NUM_NEIGHBOR_CELLS+1)+5] | arbitration_result[23*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[281] = arbitration_result[25*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[27*(NUM_NEIGHBOR_CELLS+1)+11];
assign force_cache_write_success[282] = arbitration_result[60*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[47*(NUM_NEIGHBOR_CELLS+1)+6];
assign force_cache_write_success[283] = arbitration_result[39*(NUM_NEIGHBOR_CELLS+1)+7] | arbitration_result[28*(NUM_NEIGHBOR_CELLS+1)+10];
assign force_cache_write_success[284] = arbitration_result[31*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[56*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[285] = arbitration_result[63*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[36*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[286] = arbitration_result[55*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[41*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[287] = arbitration_result[41*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[20*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[288] = arbitration_result[26*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[24*(NUM_NEIGHBOR_CELLS+1)+11];
assign force_cache_write_success[289] = arbitration_result[61*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[44*(NUM_NEIGHBOR_CELLS+1)+6];
assign force_cache_write_success[290] = arbitration_result[36*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[29*(NUM_NEIGHBOR_CELLS+1)+10];
assign force_cache_write_success[291] = arbitration_result[28*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[57*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[292] = arbitration_result[60*(NUM_NEIGHBOR_CELLS+1)+7] | arbitration_result[37*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[293] = arbitration_result[52*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[42*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[294] = arbitration_result[42*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[21*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[295] = arbitration_result[27*(NUM_NEIGHBOR_CELLS+1)+12] | arbitration_result[25*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[296] = arbitration_result[62*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[45*(NUM_NEIGHBOR_CELLS+1)+6];
assign force_cache_write_success[297] = arbitration_result[37*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[30*(NUM_NEIGHBOR_CELLS+1)+10];
assign force_cache_write_success[298] = arbitration_result[29*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[58*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[299] = arbitration_result[61*(NUM_NEIGHBOR_CELLS+1)+7] | arbitration_result[38*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[300] = arbitration_result[53*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[43*(NUM_NEIGHBOR_CELLS+1)+5];
assign force_cache_write_success[301] = arbitration_result[43*(NUM_NEIGHBOR_CELLS+1)+6] | arbitration_result[22*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[302] = arbitration_result[24*(NUM_NEIGHBOR_CELLS+1)+12] | arbitration_result[26*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[303] = arbitration_result[63*(NUM_NEIGHBOR_CELLS+1)+7] | arbitration_result[46*(NUM_NEIGHBOR_CELLS+1)+6];
assign force_cache_write_success[304] = arbitration_result[38*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[31*(NUM_NEIGHBOR_CELLS+1)+11];
assign force_cache_write_success[305] = arbitration_result[30*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[59*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[306] = arbitration_result[62*(NUM_NEIGHBOR_CELLS+1)+7] | arbitration_result[39*(NUM_NEIGHBOR_CELLS+1)+8];
assign force_cache_write_success[307] = arbitration_result[54*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[40*(NUM_NEIGHBOR_CELLS+1)+6];
assign force_cache_write_success[308] = arbitration_result[44*(NUM_NEIGHBOR_CELLS+1)+7] | arbitration_result[27*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[309] = arbitration_result[29*(NUM_NEIGHBOR_CELLS+1)+12] | arbitration_result[31*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[310] = arbitration_result[48*(NUM_NEIGHBOR_CELLS+1)+7] | arbitration_result[35*(NUM_NEIGHBOR_CELLS+1)+8];
assign force_cache_write_success[311] = arbitration_result[43*(NUM_NEIGHBOR_CELLS+1)+7] | arbitration_result[16*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[312] = arbitration_result[19*(NUM_NEIGHBOR_CELLS+1)+12] | arbitration_result[60*(NUM_NEIGHBOR_CELLS+1)+8];
assign force_cache_write_success[313] = arbitration_result[51*(NUM_NEIGHBOR_CELLS+1)+7] | arbitration_result[40*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[314] = arbitration_result[59*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[45*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[315] = arbitration_result[45*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[24*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[316] = arbitration_result[30*(NUM_NEIGHBOR_CELLS+1)+12] | arbitration_result[28*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[317] = arbitration_result[49*(NUM_NEIGHBOR_CELLS+1)+7] | arbitration_result[32*(NUM_NEIGHBOR_CELLS+1)+8];
assign force_cache_write_success[318] = arbitration_result[40*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[17*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[319] = arbitration_result[16*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[61*(NUM_NEIGHBOR_CELLS+1)+8];
assign force_cache_write_success[320] = arbitration_result[48*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[41*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[321] = arbitration_result[56*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[46*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[322] = arbitration_result[46*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[25*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[323] = arbitration_result[31*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[29*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[324] = arbitration_result[50*(NUM_NEIGHBOR_CELLS+1)+7] | arbitration_result[33*(NUM_NEIGHBOR_CELLS+1)+8];
assign force_cache_write_success[325] = arbitration_result[41*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[18*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[326] = arbitration_result[17*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[62*(NUM_NEIGHBOR_CELLS+1)+8];
assign force_cache_write_success[327] = arbitration_result[49*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[42*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[328] = arbitration_result[57*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[47*(NUM_NEIGHBOR_CELLS+1)+7];
assign force_cache_write_success[329] = arbitration_result[47*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[26*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[330] = arbitration_result[28*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[30*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[331] = arbitration_result[51*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[34*(NUM_NEIGHBOR_CELLS+1)+8];
assign force_cache_write_success[332] = arbitration_result[42*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[19*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[333] = arbitration_result[18*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[63*(NUM_NEIGHBOR_CELLS+1)+8];
assign force_cache_write_success[334] = arbitration_result[50*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[43*(NUM_NEIGHBOR_CELLS+1)+8];
assign force_cache_write_success[335] = arbitration_result[58*(NUM_NEIGHBOR_CELLS+1)+8] | arbitration_result[44*(NUM_NEIGHBOR_CELLS+1)+8];
assign force_cache_write_success[336] = arbitration_result[48*(NUM_NEIGHBOR_CELLS+1)+9] | arbitration_result[47*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[337] = arbitration_result[33*(NUM_NEIGHBOR_CELLS+1)+9] | arbitration_result[35*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[338] = arbitration_result[4*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[55*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[339] = arbitration_result[63*(NUM_NEIGHBOR_CELLS+1)+9] | arbitration_result[36*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[340] = arbitration_result[39*(NUM_NEIGHBOR_CELLS+1)+9] | arbitration_result[0*(NUM_NEIGHBOR_CELLS+1)+10];
assign force_cache_write_success[341] = arbitration_result[7*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[60*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[342] = arbitration_result[15*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[49*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[343] = arbitration_result[49*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[44*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[344] = arbitration_result[34*(NUM_NEIGHBOR_CELLS+1)+9] | arbitration_result[32*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[345] = arbitration_result[5*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[52*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[346] = arbitration_result[60*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[37*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[347] = arbitration_result[36*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[1*(NUM_NEIGHBOR_CELLS+1)+10];
assign force_cache_write_success[348] = arbitration_result[4*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[61*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[349] = arbitration_result[12*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[50*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[350] = arbitration_result[50*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[45*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[351] = arbitration_result[35*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[33*(NUM_NEIGHBOR_CELLS+1)+10];
assign force_cache_write_success[352] = arbitration_result[6*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[53*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[353] = arbitration_result[61*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[38*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[354] = arbitration_result[37*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[2*(NUM_NEIGHBOR_CELLS+1)+10];
assign force_cache_write_success[355] = arbitration_result[5*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[62*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[356] = arbitration_result[13*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[51*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[357] = arbitration_result[51*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[46*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[358] = arbitration_result[32*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[34*(NUM_NEIGHBOR_CELLS+1)+10];
assign force_cache_write_success[359] = arbitration_result[7*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[54*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[360] = arbitration_result[62*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[39*(NUM_NEIGHBOR_CELLS+1)+10];
assign force_cache_write_success[361] = arbitration_result[38*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[3*(NUM_NEIGHBOR_CELLS+1)+10];
assign force_cache_write_success[362] = arbitration_result[6*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[63*(NUM_NEIGHBOR_CELLS+1)+10];
assign force_cache_write_success[363] = arbitration_result[14*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[48*(NUM_NEIGHBOR_CELLS+1)+10];
assign force_cache_write_success[364] = arbitration_result[52*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[35*(NUM_NEIGHBOR_CELLS+1)+11];
assign force_cache_write_success[365] = arbitration_result[37*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[39*(NUM_NEIGHBOR_CELLS+1)+11];
assign force_cache_write_success[366] = arbitration_result[8*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[59*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[367] = arbitration_result[51*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[40*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[368] = arbitration_result[43*(NUM_NEIGHBOR_CELLS+1)+9] | arbitration_result[4*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[369] = arbitration_result[11*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[48*(NUM_NEIGHBOR_CELLS+1)+11];
assign force_cache_write_success[370] = arbitration_result[3*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[53*(NUM_NEIGHBOR_CELLS+1)+10];
assign force_cache_write_success[371] = arbitration_result[53*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[32*(NUM_NEIGHBOR_CELLS+1)+11];
assign force_cache_write_success[372] = arbitration_result[38*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[36*(NUM_NEIGHBOR_CELLS+1)+11];
assign force_cache_write_success[373] = arbitration_result[9*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[56*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[374] = arbitration_result[48*(NUM_NEIGHBOR_CELLS+1)+12] | arbitration_result[41*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[375] = arbitration_result[40*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[5*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[376] = arbitration_result[8*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[49*(NUM_NEIGHBOR_CELLS+1)+11];
assign force_cache_write_success[377] = arbitration_result[0*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[54*(NUM_NEIGHBOR_CELLS+1)+10];
assign force_cache_write_success[378] = arbitration_result[54*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[33*(NUM_NEIGHBOR_CELLS+1)+11];
assign force_cache_write_success[379] = arbitration_result[39*(NUM_NEIGHBOR_CELLS+1)+12] | arbitration_result[37*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[380] = arbitration_result[10*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[57*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[381] = arbitration_result[49*(NUM_NEIGHBOR_CELLS+1)+12] | arbitration_result[42*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[382] = arbitration_result[41*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[6*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[383] = arbitration_result[9*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[50*(NUM_NEIGHBOR_CELLS+1)+11];
assign force_cache_write_success[384] = arbitration_result[1*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[55*(NUM_NEIGHBOR_CELLS+1)+10];
assign force_cache_write_success[385] = arbitration_result[55*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[34*(NUM_NEIGHBOR_CELLS+1)+11];
assign force_cache_write_success[386] = arbitration_result[36*(NUM_NEIGHBOR_CELLS+1)+12] | arbitration_result[38*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[387] = arbitration_result[11*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[58*(NUM_NEIGHBOR_CELLS+1)+9];
assign force_cache_write_success[388] = arbitration_result[50*(NUM_NEIGHBOR_CELLS+1)+12] | arbitration_result[43*(NUM_NEIGHBOR_CELLS+1)+10];
assign force_cache_write_success[389] = arbitration_result[42*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[7*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[390] = arbitration_result[10*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[51*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[391] = arbitration_result[2*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[52*(NUM_NEIGHBOR_CELLS+1)+11];
assign force_cache_write_success[392] = arbitration_result[56*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[39*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[393] = arbitration_result[41*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[43*(NUM_NEIGHBOR_CELLS+1)+11];
assign force_cache_write_success[394] = arbitration_result[12*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[63*(NUM_NEIGHBOR_CELLS+1)+11];
assign force_cache_write_success[395] = arbitration_result[55*(NUM_NEIGHBOR_CELLS+1)+12] | arbitration_result[44*(NUM_NEIGHBOR_CELLS+1)+10];
assign force_cache_write_success[396] = arbitration_result[47*(NUM_NEIGHBOR_CELLS+1)+10] | arbitration_result[8*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[397] = arbitration_result[15*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[52*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[398] = arbitration_result[7*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[57*(NUM_NEIGHBOR_CELLS+1)+10];
assign force_cache_write_success[399] = arbitration_result[57*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[36*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[400] = arbitration_result[42*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[40*(NUM_NEIGHBOR_CELLS+1)+11];
assign force_cache_write_success[401] = arbitration_result[13*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[60*(NUM_NEIGHBOR_CELLS+1)+11];
assign force_cache_write_success[402] = arbitration_result[52*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[45*(NUM_NEIGHBOR_CELLS+1)+10];
assign force_cache_write_success[403] = arbitration_result[44*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[9*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[404] = arbitration_result[12*(NUM_NEIGHBOR_CELLS+1)+12] | arbitration_result[53*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[405] = arbitration_result[4*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[58*(NUM_NEIGHBOR_CELLS+1)+10];
assign force_cache_write_success[406] = arbitration_result[58*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[37*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[407] = arbitration_result[43*(NUM_NEIGHBOR_CELLS+1)+12] | arbitration_result[41*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[408] = arbitration_result[14*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[61*(NUM_NEIGHBOR_CELLS+1)+11];
assign force_cache_write_success[409] = arbitration_result[53*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[46*(NUM_NEIGHBOR_CELLS+1)+10];
assign force_cache_write_success[410] = arbitration_result[45*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[10*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[411] = arbitration_result[13*(NUM_NEIGHBOR_CELLS+1)+12] | arbitration_result[54*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[412] = arbitration_result[5*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[59*(NUM_NEIGHBOR_CELLS+1)+10];
assign force_cache_write_success[413] = arbitration_result[59*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[38*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[414] = arbitration_result[40*(NUM_NEIGHBOR_CELLS+1)+12] | arbitration_result[42*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[415] = arbitration_result[15*(NUM_NEIGHBOR_CELLS+1)+12] | arbitration_result[62*(NUM_NEIGHBOR_CELLS+1)+11];
assign force_cache_write_success[416] = arbitration_result[54*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[47*(NUM_NEIGHBOR_CELLS+1)+11];
assign force_cache_write_success[417] = arbitration_result[46*(NUM_NEIGHBOR_CELLS+1)+11] | arbitration_result[11*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[418] = arbitration_result[14*(NUM_NEIGHBOR_CELLS+1)+12] | arbitration_result[55*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[419] = arbitration_result[6*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[56*(NUM_NEIGHBOR_CELLS+1)+11];
assign force_cache_write_success[420] = arbitration_result[60*(NUM_NEIGHBOR_CELLS+1)+12] | arbitration_result[43*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[421] = arbitration_result[45*(NUM_NEIGHBOR_CELLS+1)+12] | arbitration_result[47*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[422] = arbitration_result[0*(NUM_NEIGHBOR_CELLS+1)+12] | arbitration_result[51*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[423] = arbitration_result[59*(NUM_NEIGHBOR_CELLS+1)+12] | arbitration_result[32*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[424] = arbitration_result[35*(NUM_NEIGHBOR_CELLS+1)+12] | arbitration_result[12*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[425] = arbitration_result[3*(NUM_NEIGHBOR_CELLS+1)+12] | arbitration_result[56*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[426] = arbitration_result[11*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[61*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[427] = arbitration_result[61*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[40*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[428] = arbitration_result[46*(NUM_NEIGHBOR_CELLS+1)+12] | arbitration_result[44*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[429] = arbitration_result[1*(NUM_NEIGHBOR_CELLS+1)+12] | arbitration_result[48*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[430] = arbitration_result[56*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[33*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[431] = arbitration_result[32*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[13*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[432] = arbitration_result[0*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[57*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[433] = arbitration_result[8*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[62*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[434] = arbitration_result[62*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[41*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[435] = arbitration_result[47*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[45*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[436] = arbitration_result[2*(NUM_NEIGHBOR_CELLS+1)+12] | arbitration_result[49*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[437] = arbitration_result[57*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[34*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[438] = arbitration_result[33*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[14*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[439] = arbitration_result[1*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[58*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[440] = arbitration_result[9*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[63*(NUM_NEIGHBOR_CELLS+1)+12];
assign force_cache_write_success[441] = arbitration_result[63*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[42*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[442] = arbitration_result[44*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[46*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[443] = arbitration_result[3*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[50*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[444] = arbitration_result[58*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[35*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[445] = arbitration_result[34*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[15*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[446] = arbitration_result[2*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[59*(NUM_NEIGHBOR_CELLS+1)+13];
assign force_cache_write_success[447] = arbitration_result[10*(NUM_NEIGHBOR_CELLS+1)+13] | arbitration_result[60*(NUM_NEIGHBOR_CELLS+1)+13];

endmodule