// DualPort_RAM_Test.v

// Generated using ACDS version 18.0 219

`timescale 1 ps / 1 ps
module DualPort_RAM_Test (
		input  wire [95:0] data,      //  ram_input.datain
		input  wire [8:0]  wraddress, //           .wraddress
		input  wire [8:0]  rdaddress, //           .rdaddress
		input  wire        wren,      //           .wren
		input  wire        clock,     //           .clock
		output wire [95:0] q          // ram_output.dataout
	);

	DualPort_RAM_Test_ram_2port_180_bi2xvuy ram_2port_0 (
		.data      (data),      //   input,  width = 96,  ram_input.datain
		.wraddress (wraddress), //   input,   width = 9,           .wraddress
		.rdaddress (rdaddress), //   input,   width = 9,           .rdaddress
		.wren      (wren),      //   input,   width = 1,           .wren
		.clock     (clock),     //   input,   width = 1,           .clock
		.q         (q)          //  output,  width = 96, ram_output.dataout
	);

endmodule
