module Int_Mul_Add (
		input  wire [3:0] dataa_0, // dataa_0.dataa_0
		input  wire [3:0] datab_0, // datab_0.datab_0
		output wire [3:0] result   //  result.result
	);
endmodule

