// FP_Sqrt.v

// Generated using ACDS version 18.0 219

`timescale 1 ps / 1 ps
module FP_Sqrt (
		input  wire [31:0] a,      //      a.a
		input  wire        areset, // areset.reset
		input  wire        clk,    //    clk.clk
		output wire [31:0] q       //      q.q
	);

	FP_Sqrt_altera_fp_functions_180_vxsqyia fp_functions_0 (
		.clk    (clk),    //   input,   width = 1,    clk.clk
		.areset (areset), //   input,   width = 1, areset.reset
		.a      (a),      //   input,  width = 32,      a.a
		.q      (q)       //  output,  width = 32,      q.q
	);

endmodule
