module force_valid_to_enable_mapping
#(
	parameter NUM_CELLS = 64, 
	parameter NUM_NEIGHBOR_CELLS = 13, 
	parameter NUM_FILTER = 7
)
(
	input [NUM_CELLS*NUM_FILTER-1:0] force_valid, 
	input [NUM_CELLS*NUM_FILTER-1:0] force_dst, 
	
	output [NUM_CELLS*(NUM_NEIGHBOR_CELLS+1)-1:0] force_wr_enable_splitted
);

assign force_wr_enable_splitted[0*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[0]) ? 1'b0 : force_valid[0];
assign force_wr_enable_splitted[0*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[27]) ? force_valid[27] : 1'b0;
assign force_wr_enable_splitted[0*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[33]) ? force_valid[33] : 1'b0;
assign force_wr_enable_splitted[0*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[38]) ? 1'b0 : force_valid[38];
assign force_wr_enable_splitted[0*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[93]) ? force_valid[93] : 1'b0;
assign force_wr_enable_splitted[0*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[120]) ? force_valid[120] : 1'b0;
assign force_wr_enable_splitted[0*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[134]) ? 1'b0 : force_valid[134];
assign force_wr_enable_splitted[0*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[147]) ? force_valid[147] : 1'b0;
assign force_wr_enable_splitted[0*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[199]) ? force_valid[199] : 1'b0;
assign force_wr_enable_splitted[0*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[207]) ? 1'b0 : force_valid[207];
assign force_wr_enable_splitted[0*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[340]) ? force_valid[340] : 1'b0;
assign force_wr_enable_splitted[0*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[377]) ? 1'b0 : force_valid[377];
assign force_wr_enable_splitted[0*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[422]) ? 1'b0 : force_valid[422];
assign force_wr_enable_splitted[0*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[432]) ? 1'b0 : force_valid[432];
assign force_wr_enable_splitted[1*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[6]) ? force_valid[6] : 1'b0;
assign force_wr_enable_splitted[1*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[7]) ? 1'b0 : force_valid[7];
assign force_wr_enable_splitted[1*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[40]) ? force_valid[40] : 1'b0;
assign force_wr_enable_splitted[1*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[45]) ? 1'b0 : force_valid[45];
assign force_wr_enable_splitted[1*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[100]) ? force_valid[100] : 1'b0;
assign force_wr_enable_splitted[1*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[113]) ? 1'b0 : force_valid[113];
assign force_wr_enable_splitted[1*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[127]) ? force_valid[127] : 1'b0;
assign force_wr_enable_splitted[1*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[154]) ? force_valid[154] : 1'b0;
assign force_wr_enable_splitted[1*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[206]) ? force_valid[206] : 1'b0;
assign force_wr_enable_splitted[1*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[214]) ? 1'b0 : force_valid[214];
assign force_wr_enable_splitted[1*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[347]) ? force_valid[347] : 1'b0;
assign force_wr_enable_splitted[1*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[384]) ? 1'b0 : force_valid[384];
assign force_wr_enable_splitted[1*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[429]) ? 1'b0 : force_valid[429];
assign force_wr_enable_splitted[1*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[439]) ? 1'b0 : force_valid[439];
assign force_wr_enable_splitted[2*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[13]) ? force_valid[13] : 1'b0;
assign force_wr_enable_splitted[2*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[14]) ? 1'b0 : force_valid[14];
assign force_wr_enable_splitted[2*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[47]) ? force_valid[47] : 1'b0;
assign force_wr_enable_splitted[2*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[52]) ? 1'b0 : force_valid[52];
assign force_wr_enable_splitted[2*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[107]) ? force_valid[107] : 1'b0;
assign force_wr_enable_splitted[2*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[120]) ? 1'b0 : force_valid[120];
assign force_wr_enable_splitted[2*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[134]) ? force_valid[134] : 1'b0;
assign force_wr_enable_splitted[2*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[161]) ? force_valid[161] : 1'b0;
assign force_wr_enable_splitted[2*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[213]) ? force_valid[213] : 1'b0;
assign force_wr_enable_splitted[2*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[221]) ? 1'b0 : force_valid[221];
assign force_wr_enable_splitted[2*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[354]) ? force_valid[354] : 1'b0;
assign force_wr_enable_splitted[2*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[391]) ? 1'b0 : force_valid[391];
assign force_wr_enable_splitted[2*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[436]) ? 1'b0 : force_valid[436];
assign force_wr_enable_splitted[2*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[446]) ? 1'b0 : force_valid[446];
assign force_wr_enable_splitted[3*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[20]) ? force_valid[20] : 1'b0;
assign force_wr_enable_splitted[3*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[21]) ? 1'b0 : force_valid[21];
assign force_wr_enable_splitted[3*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[31]) ? 1'b0 : force_valid[31];
assign force_wr_enable_splitted[3*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[54]) ? force_valid[54] : 1'b0;
assign force_wr_enable_splitted[3*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[86]) ? force_valid[86] : 1'b0;
assign force_wr_enable_splitted[3*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[113]) ? force_valid[113] : 1'b0;
assign force_wr_enable_splitted[3*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[127]) ? 1'b0 : force_valid[127];
assign force_wr_enable_splitted[3*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[140]) ? force_valid[140] : 1'b0;
assign force_wr_enable_splitted[3*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[200]) ? 1'b0 : force_valid[200];
assign force_wr_enable_splitted[3*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[220]) ? force_valid[220] : 1'b0;
assign force_wr_enable_splitted[3*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[361]) ? force_valid[361] : 1'b0;
assign force_wr_enable_splitted[3*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[370]) ? 1'b0 : force_valid[370];
assign force_wr_enable_splitted[3*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[425]) ? 1'b0 : force_valid[425];
assign force_wr_enable_splitted[3*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[443]) ? 1'b0 : force_valid[443];
assign force_wr_enable_splitted[4*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[9]) ? force_valid[9] : 1'b0;
assign force_wr_enable_splitted[4*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[28]) ? 1'b0 : force_valid[28];
assign force_wr_enable_splitted[4*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[55]) ? force_valid[55] : 1'b0;
assign force_wr_enable_splitted[4*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[61]) ? force_valid[61] : 1'b0;
assign force_wr_enable_splitted[4*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[66]) ? 1'b0 : force_valid[66];
assign force_wr_enable_splitted[4*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[115]) ? force_valid[115] : 1'b0;
assign force_wr_enable_splitted[4*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[123]) ? 1'b0 : force_valid[123];
assign force_wr_enable_splitted[4*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[148]) ? force_valid[148] : 1'b0;
assign force_wr_enable_splitted[4*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[162]) ? 1'b0 : force_valid[162];
assign force_wr_enable_splitted[4*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[175]) ? force_valid[175] : 1'b0;
assign force_wr_enable_splitted[4*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[338]) ? 1'b0 : force_valid[338];
assign force_wr_enable_splitted[4*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[348]) ? 1'b0 : force_valid[348];
assign force_wr_enable_splitted[4*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[368]) ? force_valid[368] : 1'b0;
assign force_wr_enable_splitted[4*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[405]) ? 1'b0 : force_valid[405];
assign force_wr_enable_splitted[5*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[16]) ? force_valid[16] : 1'b0;
assign force_wr_enable_splitted[5*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[34]) ? force_valid[34] : 1'b0;
assign force_wr_enable_splitted[5*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[35]) ? 1'b0 : force_valid[35];
assign force_wr_enable_splitted[5*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[68]) ? force_valid[68] : 1'b0;
assign force_wr_enable_splitted[5*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[73]) ? 1'b0 : force_valid[73];
assign force_wr_enable_splitted[5*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[122]) ? force_valid[122] : 1'b0;
assign force_wr_enable_splitted[5*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[130]) ? 1'b0 : force_valid[130];
assign force_wr_enable_splitted[5*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[141]) ? 1'b0 : force_valid[141];
assign force_wr_enable_splitted[5*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[155]) ? force_valid[155] : 1'b0;
assign force_wr_enable_splitted[5*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[182]) ? force_valid[182] : 1'b0;
assign force_wr_enable_splitted[5*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[345]) ? 1'b0 : force_valid[345];
assign force_wr_enable_splitted[5*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[355]) ? 1'b0 : force_valid[355];
assign force_wr_enable_splitted[5*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[375]) ? force_valid[375] : 1'b0;
assign force_wr_enable_splitted[5*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[412]) ? 1'b0 : force_valid[412];
assign force_wr_enable_splitted[6*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[23]) ? force_valid[23] : 1'b0;
assign force_wr_enable_splitted[6*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[41]) ? force_valid[41] : 1'b0;
assign force_wr_enable_splitted[6*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[42]) ? 1'b0 : force_valid[42];
assign force_wr_enable_splitted[6*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[75]) ? force_valid[75] : 1'b0;
assign force_wr_enable_splitted[6*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[80]) ? 1'b0 : force_valid[80];
assign force_wr_enable_splitted[6*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[129]) ? force_valid[129] : 1'b0;
assign force_wr_enable_splitted[6*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[137]) ? 1'b0 : force_valid[137];
assign force_wr_enable_splitted[6*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[148]) ? 1'b0 : force_valid[148];
assign force_wr_enable_splitted[6*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[162]) ? force_valid[162] : 1'b0;
assign force_wr_enable_splitted[6*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[189]) ? force_valid[189] : 1'b0;
assign force_wr_enable_splitted[6*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[352]) ? 1'b0 : force_valid[352];
assign force_wr_enable_splitted[6*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[362]) ? 1'b0 : force_valid[362];
assign force_wr_enable_splitted[6*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[382]) ? force_valid[382] : 1'b0;
assign force_wr_enable_splitted[6*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[419]) ? 1'b0 : force_valid[419];
assign force_wr_enable_splitted[7*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[2]) ? force_valid[2] : 1'b0;
assign force_wr_enable_splitted[7*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[48]) ? force_valid[48] : 1'b0;
assign force_wr_enable_splitted[7*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[49]) ? 1'b0 : force_valid[49];
assign force_wr_enable_splitted[7*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[59]) ? 1'b0 : force_valid[59];
assign force_wr_enable_splitted[7*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[82]) ? force_valid[82] : 1'b0;
assign force_wr_enable_splitted[7*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[116]) ? 1'b0 : force_valid[116];
assign force_wr_enable_splitted[7*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[136]) ? force_valid[136] : 1'b0;
assign force_wr_enable_splitted[7*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[141]) ? force_valid[141] : 1'b0;
assign force_wr_enable_splitted[7*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[155]) ? 1'b0 : force_valid[155];
assign force_wr_enable_splitted[7*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[168]) ? force_valid[168] : 1'b0;
assign force_wr_enable_splitted[7*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[341]) ? 1'b0 : force_valid[341];
assign force_wr_enable_splitted[7*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[359]) ? 1'b0 : force_valid[359];
assign force_wr_enable_splitted[7*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[389]) ? force_valid[389] : 1'b0;
assign force_wr_enable_splitted[7*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[398]) ? 1'b0 : force_valid[398];
assign force_wr_enable_splitted[8*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[37]) ? force_valid[37] : 1'b0;
assign force_wr_enable_splitted[8*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[56]) ? 1'b0 : force_valid[56];
assign force_wr_enable_splitted[8*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[83]) ? force_valid[83] : 1'b0;
assign force_wr_enable_splitted[8*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[89]) ? force_valid[89] : 1'b0;
assign force_wr_enable_splitted[8*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[94]) ? 1'b0 : force_valid[94];
assign force_wr_enable_splitted[8*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[143]) ? force_valid[143] : 1'b0;
assign force_wr_enable_splitted[8*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[151]) ? 1'b0 : force_valid[151];
assign force_wr_enable_splitted[8*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[176]) ? force_valid[176] : 1'b0;
assign force_wr_enable_splitted[8*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[190]) ? 1'b0 : force_valid[190];
assign force_wr_enable_splitted[8*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[203]) ? force_valid[203] : 1'b0;
assign force_wr_enable_splitted[8*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[366]) ? 1'b0 : force_valid[366];
assign force_wr_enable_splitted[8*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[376]) ? 1'b0 : force_valid[376];
assign force_wr_enable_splitted[8*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[396]) ? force_valid[396] : 1'b0;
assign force_wr_enable_splitted[8*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[433]) ? 1'b0 : force_valid[433];
assign force_wr_enable_splitted[9*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[44]) ? force_valid[44] : 1'b0;
assign force_wr_enable_splitted[9*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[62]) ? force_valid[62] : 1'b0;
assign force_wr_enable_splitted[9*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[63]) ? 1'b0 : force_valid[63];
assign force_wr_enable_splitted[9*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[96]) ? force_valid[96] : 1'b0;
assign force_wr_enable_splitted[9*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[101]) ? 1'b0 : force_valid[101];
assign force_wr_enable_splitted[9*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[150]) ? force_valid[150] : 1'b0;
assign force_wr_enable_splitted[9*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[158]) ? 1'b0 : force_valid[158];
assign force_wr_enable_splitted[9*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[169]) ? 1'b0 : force_valid[169];
assign force_wr_enable_splitted[9*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[183]) ? force_valid[183] : 1'b0;
assign force_wr_enable_splitted[9*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[210]) ? force_valid[210] : 1'b0;
assign force_wr_enable_splitted[9*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[373]) ? 1'b0 : force_valid[373];
assign force_wr_enable_splitted[9*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[383]) ? 1'b0 : force_valid[383];
assign force_wr_enable_splitted[9*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[403]) ? force_valid[403] : 1'b0;
assign force_wr_enable_splitted[9*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[440]) ? 1'b0 : force_valid[440];
assign force_wr_enable_splitted[10*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[51]) ? force_valid[51] : 1'b0;
assign force_wr_enable_splitted[10*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[69]) ? force_valid[69] : 1'b0;
assign force_wr_enable_splitted[10*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[70]) ? 1'b0 : force_valid[70];
assign force_wr_enable_splitted[10*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[103]) ? force_valid[103] : 1'b0;
assign force_wr_enable_splitted[10*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[108]) ? 1'b0 : force_valid[108];
assign force_wr_enable_splitted[10*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[157]) ? force_valid[157] : 1'b0;
assign force_wr_enable_splitted[10*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[165]) ? 1'b0 : force_valid[165];
assign force_wr_enable_splitted[10*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[176]) ? 1'b0 : force_valid[176];
assign force_wr_enable_splitted[10*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[190]) ? force_valid[190] : 1'b0;
assign force_wr_enable_splitted[10*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[217]) ? force_valid[217] : 1'b0;
assign force_wr_enable_splitted[10*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[380]) ? 1'b0 : force_valid[380];
assign force_wr_enable_splitted[10*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[390]) ? 1'b0 : force_valid[390];
assign force_wr_enable_splitted[10*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[410]) ? force_valid[410] : 1'b0;
assign force_wr_enable_splitted[10*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[447]) ? 1'b0 : force_valid[447];
assign force_wr_enable_splitted[11*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[30]) ? force_valid[30] : 1'b0;
assign force_wr_enable_splitted[11*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[76]) ? force_valid[76] : 1'b0;
assign force_wr_enable_splitted[11*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[77]) ? 1'b0 : force_valid[77];
assign force_wr_enable_splitted[11*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[87]) ? 1'b0 : force_valid[87];
assign force_wr_enable_splitted[11*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[110]) ? force_valid[110] : 1'b0;
assign force_wr_enable_splitted[11*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[144]) ? 1'b0 : force_valid[144];
assign force_wr_enable_splitted[11*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[164]) ? force_valid[164] : 1'b0;
assign force_wr_enable_splitted[11*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[169]) ? force_valid[169] : 1'b0;
assign force_wr_enable_splitted[11*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[183]) ? 1'b0 : force_valid[183];
assign force_wr_enable_splitted[11*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[196]) ? force_valid[196] : 1'b0;
assign force_wr_enable_splitted[11*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[369]) ? 1'b0 : force_valid[369];
assign force_wr_enable_splitted[11*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[387]) ? 1'b0 : force_valid[387];
assign force_wr_enable_splitted[11*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[417]) ? force_valid[417] : 1'b0;
assign force_wr_enable_splitted[11*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[426]) ? 1'b0 : force_valid[426];
assign force_wr_enable_splitted[12*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[5]) ? force_valid[5] : 1'b0;
assign force_wr_enable_splitted[12*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[10]) ? 1'b0 : force_valid[10];
assign force_wr_enable_splitted[12*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[65]) ? force_valid[65] : 1'b0;
assign force_wr_enable_splitted[12*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[84]) ? 1'b0 : force_valid[84];
assign force_wr_enable_splitted[12*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[111]) ? force_valid[111] : 1'b0;
assign force_wr_enable_splitted[12*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[119]) ? force_valid[119] : 1'b0;
assign force_wr_enable_splitted[12*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[171]) ? force_valid[171] : 1'b0;
assign force_wr_enable_splitted[12*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[179]) ? 1'b0 : force_valid[179];
assign force_wr_enable_splitted[12*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[204]) ? force_valid[204] : 1'b0;
assign force_wr_enable_splitted[12*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[218]) ? 1'b0 : force_valid[218];
assign force_wr_enable_splitted[12*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[349]) ? 1'b0 : force_valid[349];
assign force_wr_enable_splitted[12*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[394]) ? 1'b0 : force_valid[394];
assign force_wr_enable_splitted[12*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[404]) ? 1'b0 : force_valid[404];
assign force_wr_enable_splitted[12*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[424]) ? force_valid[424] : 1'b0;
assign force_wr_enable_splitted[13*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[12]) ? force_valid[12] : 1'b0;
assign force_wr_enable_splitted[13*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[17]) ? 1'b0 : force_valid[17];
assign force_wr_enable_splitted[13*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[72]) ? force_valid[72] : 1'b0;
assign force_wr_enable_splitted[13*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[90]) ? force_valid[90] : 1'b0;
assign force_wr_enable_splitted[13*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[91]) ? 1'b0 : force_valid[91];
assign force_wr_enable_splitted[13*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[126]) ? force_valid[126] : 1'b0;
assign force_wr_enable_splitted[13*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[178]) ? force_valid[178] : 1'b0;
assign force_wr_enable_splitted[13*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[186]) ? 1'b0 : force_valid[186];
assign force_wr_enable_splitted[13*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[197]) ? 1'b0 : force_valid[197];
assign force_wr_enable_splitted[13*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[211]) ? force_valid[211] : 1'b0;
assign force_wr_enable_splitted[13*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[356]) ? 1'b0 : force_valid[356];
assign force_wr_enable_splitted[13*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[401]) ? 1'b0 : force_valid[401];
assign force_wr_enable_splitted[13*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[411]) ? 1'b0 : force_valid[411];
assign force_wr_enable_splitted[13*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[431]) ? force_valid[431] : 1'b0;
assign force_wr_enable_splitted[14*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[19]) ? force_valid[19] : 1'b0;
assign force_wr_enable_splitted[14*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[24]) ? 1'b0 : force_valid[24];
assign force_wr_enable_splitted[14*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[79]) ? force_valid[79] : 1'b0;
assign force_wr_enable_splitted[14*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[97]) ? force_valid[97] : 1'b0;
assign force_wr_enable_splitted[14*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[98]) ? 1'b0 : force_valid[98];
assign force_wr_enable_splitted[14*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[133]) ? force_valid[133] : 1'b0;
assign force_wr_enable_splitted[14*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[185]) ? force_valid[185] : 1'b0;
assign force_wr_enable_splitted[14*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[193]) ? 1'b0 : force_valid[193];
assign force_wr_enable_splitted[14*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[204]) ? 1'b0 : force_valid[204];
assign force_wr_enable_splitted[14*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[218]) ? force_valid[218] : 1'b0;
assign force_wr_enable_splitted[14*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[363]) ? 1'b0 : force_valid[363];
assign force_wr_enable_splitted[14*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[408]) ? 1'b0 : force_valid[408];
assign force_wr_enable_splitted[14*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[418]) ? 1'b0 : force_valid[418];
assign force_wr_enable_splitted[14*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[438]) ? force_valid[438] : 1'b0;
assign force_wr_enable_splitted[15*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[3]) ? 1'b0 : force_valid[3];
assign force_wr_enable_splitted[15*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[26]) ? force_valid[26] : 1'b0;
assign force_wr_enable_splitted[15*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[58]) ? force_valid[58] : 1'b0;
assign force_wr_enable_splitted[15*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[104]) ? force_valid[104] : 1'b0;
assign force_wr_enable_splitted[15*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[105]) ? 1'b0 : force_valid[105];
assign force_wr_enable_splitted[15*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[112]) ? force_valid[112] : 1'b0;
assign force_wr_enable_splitted[15*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[172]) ? 1'b0 : force_valid[172];
assign force_wr_enable_splitted[15*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[192]) ? force_valid[192] : 1'b0;
assign force_wr_enable_splitted[15*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[197]) ? force_valid[197] : 1'b0;
assign force_wr_enable_splitted[15*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[211]) ? 1'b0 : force_valid[211];
assign force_wr_enable_splitted[15*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[342]) ? 1'b0 : force_valid[342];
assign force_wr_enable_splitted[15*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[397]) ? 1'b0 : force_valid[397];
assign force_wr_enable_splitted[15*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[415]) ? 1'b0 : force_valid[415];
assign force_wr_enable_splitted[15*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[445]) ? force_valid[445] : 1'b0;
assign force_wr_enable_splitted[16*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[4]) ? force_valid[4] : 1'b0;
assign force_wr_enable_splitted[16*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[41]) ? 1'b0 : force_valid[41];
assign force_wr_enable_splitted[16*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[86]) ? 1'b0 : force_valid[86];
assign force_wr_enable_splitted[16*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[96]) ? 1'b0 : force_valid[96];
assign force_wr_enable_splitted[16*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[112]) ? 1'b0 : force_valid[112];
assign force_wr_enable_splitted[16*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[139]) ? force_valid[139] : 1'b0;
assign force_wr_enable_splitted[16*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[145]) ? force_valid[145] : 1'b0;
assign force_wr_enable_splitted[16*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[150]) ? 1'b0 : force_valid[150];
assign force_wr_enable_splitted[16*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[205]) ? force_valid[205] : 1'b0;
assign force_wr_enable_splitted[16*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[232]) ? force_valid[232] : 1'b0;
assign force_wr_enable_splitted[16*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[246]) ? 1'b0 : force_valid[246];
assign force_wr_enable_splitted[16*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[259]) ? force_valid[259] : 1'b0;
assign force_wr_enable_splitted[16*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[311]) ? force_valid[311] : 1'b0;
assign force_wr_enable_splitted[16*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[319]) ? 1'b0 : force_valid[319];
assign force_wr_enable_splitted[17*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[11]) ? force_valid[11] : 1'b0;
assign force_wr_enable_splitted[17*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[48]) ? 1'b0 : force_valid[48];
assign force_wr_enable_splitted[17*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[93]) ? 1'b0 : force_valid[93];
assign force_wr_enable_splitted[17*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[103]) ? 1'b0 : force_valid[103];
assign force_wr_enable_splitted[17*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[118]) ? force_valid[118] : 1'b0;
assign force_wr_enable_splitted[17*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[119]) ? 1'b0 : force_valid[119];
assign force_wr_enable_splitted[17*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[152]) ? force_valid[152] : 1'b0;
assign force_wr_enable_splitted[17*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[157]) ? 1'b0 : force_valid[157];
assign force_wr_enable_splitted[17*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[212]) ? force_valid[212] : 1'b0;
assign force_wr_enable_splitted[17*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[225]) ? 1'b0 : force_valid[225];
assign force_wr_enable_splitted[17*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[239]) ? force_valid[239] : 1'b0;
assign force_wr_enable_splitted[17*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[266]) ? force_valid[266] : 1'b0;
assign force_wr_enable_splitted[17*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[318]) ? force_valid[318] : 1'b0;
assign force_wr_enable_splitted[17*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[326]) ? 1'b0 : force_valid[326];
assign force_wr_enable_splitted[18*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[18]) ? force_valid[18] : 1'b0;
assign force_wr_enable_splitted[18*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[55]) ? 1'b0 : force_valid[55];
assign force_wr_enable_splitted[18*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[100]) ? 1'b0 : force_valid[100];
assign force_wr_enable_splitted[18*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[110]) ? 1'b0 : force_valid[110];
assign force_wr_enable_splitted[18*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[125]) ? force_valid[125] : 1'b0;
assign force_wr_enable_splitted[18*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[126]) ? 1'b0 : force_valid[126];
assign force_wr_enable_splitted[18*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[159]) ? force_valid[159] : 1'b0;
assign force_wr_enable_splitted[18*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[164]) ? 1'b0 : force_valid[164];
assign force_wr_enable_splitted[18*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[219]) ? force_valid[219] : 1'b0;
assign force_wr_enable_splitted[18*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[232]) ? 1'b0 : force_valid[232];
assign force_wr_enable_splitted[18*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[246]) ? force_valid[246] : 1'b0;
assign force_wr_enable_splitted[18*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[273]) ? force_valid[273] : 1'b0;
assign force_wr_enable_splitted[18*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[325]) ? force_valid[325] : 1'b0;
assign force_wr_enable_splitted[18*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[333]) ? 1'b0 : force_valid[333];
assign force_wr_enable_splitted[19*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[25]) ? force_valid[25] : 1'b0;
assign force_wr_enable_splitted[19*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[34]) ? 1'b0 : force_valid[34];
assign force_wr_enable_splitted[19*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[89]) ? 1'b0 : force_valid[89];
assign force_wr_enable_splitted[19*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[107]) ? 1'b0 : force_valid[107];
assign force_wr_enable_splitted[19*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[132]) ? force_valid[132] : 1'b0;
assign force_wr_enable_splitted[19*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[133]) ? 1'b0 : force_valid[133];
assign force_wr_enable_splitted[19*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[143]) ? 1'b0 : force_valid[143];
assign force_wr_enable_splitted[19*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[166]) ? force_valid[166] : 1'b0;
assign force_wr_enable_splitted[19*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[198]) ? force_valid[198] : 1'b0;
assign force_wr_enable_splitted[19*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[225]) ? force_valid[225] : 1'b0;
assign force_wr_enable_splitted[19*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[239]) ? 1'b0 : force_valid[239];
assign force_wr_enable_splitted[19*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[252]) ? force_valid[252] : 1'b0;
assign force_wr_enable_splitted[19*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[312]) ? 1'b0 : force_valid[312];
assign force_wr_enable_splitted[19*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[332]) ? force_valid[332] : 1'b0;
assign force_wr_enable_splitted[20*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[2]) ? 1'b0 : force_valid[2];
assign force_wr_enable_splitted[20*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[12]) ? 1'b0 : force_valid[12];
assign force_wr_enable_splitted[20*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[32]) ? force_valid[32] : 1'b0;
assign force_wr_enable_splitted[20*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[69]) ? 1'b0 : force_valid[69];
assign force_wr_enable_splitted[20*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[121]) ? force_valid[121] : 1'b0;
assign force_wr_enable_splitted[20*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[140]) ? 1'b0 : force_valid[140];
assign force_wr_enable_splitted[20*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[167]) ? force_valid[167] : 1'b0;
assign force_wr_enable_splitted[20*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[173]) ? force_valid[173] : 1'b0;
assign force_wr_enable_splitted[20*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[178]) ? 1'b0 : force_valid[178];
assign force_wr_enable_splitted[20*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[227]) ? force_valid[227] : 1'b0;
assign force_wr_enable_splitted[20*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[235]) ? 1'b0 : force_valid[235];
assign force_wr_enable_splitted[20*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[260]) ? force_valid[260] : 1'b0;
assign force_wr_enable_splitted[20*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[274]) ? 1'b0 : force_valid[274];
assign force_wr_enable_splitted[20*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[287]) ? force_valid[287] : 1'b0;
assign force_wr_enable_splitted[21*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[9]) ? 1'b0 : force_valid[9];
assign force_wr_enable_splitted[21*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[19]) ? 1'b0 : force_valid[19];
assign force_wr_enable_splitted[21*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[39]) ? force_valid[39] : 1'b0;
assign force_wr_enable_splitted[21*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[76]) ? 1'b0 : force_valid[76];
assign force_wr_enable_splitted[21*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[128]) ? force_valid[128] : 1'b0;
assign force_wr_enable_splitted[21*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[146]) ? force_valid[146] : 1'b0;
assign force_wr_enable_splitted[21*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[147]) ? 1'b0 : force_valid[147];
assign force_wr_enable_splitted[21*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[180]) ? force_valid[180] : 1'b0;
assign force_wr_enable_splitted[21*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[185]) ? 1'b0 : force_valid[185];
assign force_wr_enable_splitted[21*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[234]) ? force_valid[234] : 1'b0;
assign force_wr_enable_splitted[21*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[242]) ? 1'b0 : force_valid[242];
assign force_wr_enable_splitted[21*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[253]) ? 1'b0 : force_valid[253];
assign force_wr_enable_splitted[21*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[267]) ? force_valid[267] : 1'b0;
assign force_wr_enable_splitted[21*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[294]) ? force_valid[294] : 1'b0;
assign force_wr_enable_splitted[22*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[16]) ? 1'b0 : force_valid[16];
assign force_wr_enable_splitted[22*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[26]) ? 1'b0 : force_valid[26];
assign force_wr_enable_splitted[22*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[46]) ? force_valid[46] : 1'b0;
assign force_wr_enable_splitted[22*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[83]) ? 1'b0 : force_valid[83];
assign force_wr_enable_splitted[22*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[135]) ? force_valid[135] : 1'b0;
assign force_wr_enable_splitted[22*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[153]) ? force_valid[153] : 1'b0;
assign force_wr_enable_splitted[22*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[154]) ? 1'b0 : force_valid[154];
assign force_wr_enable_splitted[22*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[187]) ? force_valid[187] : 1'b0;
assign force_wr_enable_splitted[22*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[192]) ? 1'b0 : force_valid[192];
assign force_wr_enable_splitted[22*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[241]) ? force_valid[241] : 1'b0;
assign force_wr_enable_splitted[22*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[249]) ? 1'b0 : force_valid[249];
assign force_wr_enable_splitted[22*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[260]) ? 1'b0 : force_valid[260];
assign force_wr_enable_splitted[22*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[274]) ? force_valid[274] : 1'b0;
assign force_wr_enable_splitted[22*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[301]) ? force_valid[301] : 1'b0;
assign force_wr_enable_splitted[23*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[5]) ? 1'b0 : force_valid[5];
assign force_wr_enable_splitted[23*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[23]) ? 1'b0 : force_valid[23];
assign force_wr_enable_splitted[23*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[53]) ? force_valid[53] : 1'b0;
assign force_wr_enable_splitted[23*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[62]) ? 1'b0 : force_valid[62];
assign force_wr_enable_splitted[23*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[114]) ? force_valid[114] : 1'b0;
assign force_wr_enable_splitted[23*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[160]) ? force_valid[160] : 1'b0;
assign force_wr_enable_splitted[23*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[161]) ? 1'b0 : force_valid[161];
assign force_wr_enable_splitted[23*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[171]) ? 1'b0 : force_valid[171];
assign force_wr_enable_splitted[23*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[194]) ? force_valid[194] : 1'b0;
assign force_wr_enable_splitted[23*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[228]) ? 1'b0 : force_valid[228];
assign force_wr_enable_splitted[23*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[248]) ? force_valid[248] : 1'b0;
assign force_wr_enable_splitted[23*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[253]) ? force_valid[253] : 1'b0;
assign force_wr_enable_splitted[23*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[267]) ? 1'b0 : force_valid[267];
assign force_wr_enable_splitted[23*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[280]) ? force_valid[280] : 1'b0;
assign force_wr_enable_splitted[24*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[30]) ? 1'b0 : force_valid[30];
assign force_wr_enable_splitted[24*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[40]) ? 1'b0 : force_valid[40];
assign force_wr_enable_splitted[24*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[60]) ? force_valid[60] : 1'b0;
assign force_wr_enable_splitted[24*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[97]) ? 1'b0 : force_valid[97];
assign force_wr_enable_splitted[24*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[149]) ? force_valid[149] : 1'b0;
assign force_wr_enable_splitted[24*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[168]) ? 1'b0 : force_valid[168];
assign force_wr_enable_splitted[24*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[195]) ? force_valid[195] : 1'b0;
assign force_wr_enable_splitted[24*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[201]) ? force_valid[201] : 1'b0;
assign force_wr_enable_splitted[24*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[206]) ? 1'b0 : force_valid[206];
assign force_wr_enable_splitted[24*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[255]) ? force_valid[255] : 1'b0;
assign force_wr_enable_splitted[24*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[263]) ? 1'b0 : force_valid[263];
assign force_wr_enable_splitted[24*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[288]) ? force_valid[288] : 1'b0;
assign force_wr_enable_splitted[24*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[302]) ? 1'b0 : force_valid[302];
assign force_wr_enable_splitted[24*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[315]) ? force_valid[315] : 1'b0;
assign force_wr_enable_splitted[25*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[37]) ? 1'b0 : force_valid[37];
assign force_wr_enable_splitted[25*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[47]) ? 1'b0 : force_valid[47];
assign force_wr_enable_splitted[25*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[67]) ? force_valid[67] : 1'b0;
assign force_wr_enable_splitted[25*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[104]) ? 1'b0 : force_valid[104];
assign force_wr_enable_splitted[25*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[156]) ? force_valid[156] : 1'b0;
assign force_wr_enable_splitted[25*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[174]) ? force_valid[174] : 1'b0;
assign force_wr_enable_splitted[25*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[175]) ? 1'b0 : force_valid[175];
assign force_wr_enable_splitted[25*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[208]) ? force_valid[208] : 1'b0;
assign force_wr_enable_splitted[25*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[213]) ? 1'b0 : force_valid[213];
assign force_wr_enable_splitted[25*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[262]) ? force_valid[262] : 1'b0;
assign force_wr_enable_splitted[25*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[270]) ? 1'b0 : force_valid[270];
assign force_wr_enable_splitted[25*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[281]) ? 1'b0 : force_valid[281];
assign force_wr_enable_splitted[25*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[295]) ? force_valid[295] : 1'b0;
assign force_wr_enable_splitted[25*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[322]) ? force_valid[322] : 1'b0;
assign force_wr_enable_splitted[26*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[44]) ? 1'b0 : force_valid[44];
assign force_wr_enable_splitted[26*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[54]) ? 1'b0 : force_valid[54];
assign force_wr_enable_splitted[26*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[74]) ? force_valid[74] : 1'b0;
assign force_wr_enable_splitted[26*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[111]) ? 1'b0 : force_valid[111];
assign force_wr_enable_splitted[26*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[163]) ? force_valid[163] : 1'b0;
assign force_wr_enable_splitted[26*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[181]) ? force_valid[181] : 1'b0;
assign force_wr_enable_splitted[26*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[182]) ? 1'b0 : force_valid[182];
assign force_wr_enable_splitted[26*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[215]) ? force_valid[215] : 1'b0;
assign force_wr_enable_splitted[26*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[220]) ? 1'b0 : force_valid[220];
assign force_wr_enable_splitted[26*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[269]) ? force_valid[269] : 1'b0;
assign force_wr_enable_splitted[26*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[277]) ? 1'b0 : force_valid[277];
assign force_wr_enable_splitted[26*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[288]) ? 1'b0 : force_valid[288];
assign force_wr_enable_splitted[26*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[302]) ? force_valid[302] : 1'b0;
assign force_wr_enable_splitted[26*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[329]) ? force_valid[329] : 1'b0;
assign force_wr_enable_splitted[27*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[33]) ? 1'b0 : force_valid[33];
assign force_wr_enable_splitted[27*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[51]) ? 1'b0 : force_valid[51];
assign force_wr_enable_splitted[27*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[81]) ? force_valid[81] : 1'b0;
assign force_wr_enable_splitted[27*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[90]) ? 1'b0 : force_valid[90];
assign force_wr_enable_splitted[27*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[142]) ? force_valid[142] : 1'b0;
assign force_wr_enable_splitted[27*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[188]) ? force_valid[188] : 1'b0;
assign force_wr_enable_splitted[27*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[189]) ? 1'b0 : force_valid[189];
assign force_wr_enable_splitted[27*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[199]) ? 1'b0 : force_valid[199];
assign force_wr_enable_splitted[27*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[222]) ? force_valid[222] : 1'b0;
assign force_wr_enable_splitted[27*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[256]) ? 1'b0 : force_valid[256];
assign force_wr_enable_splitted[27*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[276]) ? force_valid[276] : 1'b0;
assign force_wr_enable_splitted[27*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[281]) ? force_valid[281] : 1'b0;
assign force_wr_enable_splitted[27*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[295]) ? 1'b0 : force_valid[295];
assign force_wr_enable_splitted[27*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[308]) ? force_valid[308] : 1'b0;
assign force_wr_enable_splitted[28*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[13]) ? 1'b0 : force_valid[13];
assign force_wr_enable_splitted[28*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[58]) ? 1'b0 : force_valid[58];
assign force_wr_enable_splitted[28*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[68]) ? 1'b0 : force_valid[68];
assign force_wr_enable_splitted[28*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[88]) ? force_valid[88] : 1'b0;
assign force_wr_enable_splitted[28*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[117]) ? force_valid[117] : 1'b0;
assign force_wr_enable_splitted[28*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[122]) ? 1'b0 : force_valid[122];
assign force_wr_enable_splitted[28*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[177]) ? force_valid[177] : 1'b0;
assign force_wr_enable_splitted[28*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[196]) ? 1'b0 : force_valid[196];
assign force_wr_enable_splitted[28*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[223]) ? force_valid[223] : 1'b0;
assign force_wr_enable_splitted[28*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[231]) ? force_valid[231] : 1'b0;
assign force_wr_enable_splitted[28*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[283]) ? force_valid[283] : 1'b0;
assign force_wr_enable_splitted[28*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[291]) ? 1'b0 : force_valid[291];
assign force_wr_enable_splitted[28*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[316]) ? force_valid[316] : 1'b0;
assign force_wr_enable_splitted[28*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[330]) ? 1'b0 : force_valid[330];
assign force_wr_enable_splitted[29*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[20]) ? 1'b0 : force_valid[20];
assign force_wr_enable_splitted[29*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[65]) ? 1'b0 : force_valid[65];
assign force_wr_enable_splitted[29*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[75]) ? 1'b0 : force_valid[75];
assign force_wr_enable_splitted[29*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[95]) ? force_valid[95] : 1'b0;
assign force_wr_enable_splitted[29*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[124]) ? force_valid[124] : 1'b0;
assign force_wr_enable_splitted[29*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[129]) ? 1'b0 : force_valid[129];
assign force_wr_enable_splitted[29*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[184]) ? force_valid[184] : 1'b0;
assign force_wr_enable_splitted[29*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[202]) ? force_valid[202] : 1'b0;
assign force_wr_enable_splitted[29*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[203]) ? 1'b0 : force_valid[203];
assign force_wr_enable_splitted[29*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[238]) ? force_valid[238] : 1'b0;
assign force_wr_enable_splitted[29*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[290]) ? force_valid[290] : 1'b0;
assign force_wr_enable_splitted[29*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[298]) ? 1'b0 : force_valid[298];
assign force_wr_enable_splitted[29*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[309]) ? 1'b0 : force_valid[309];
assign force_wr_enable_splitted[29*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[323]) ? force_valid[323] : 1'b0;
assign force_wr_enable_splitted[30*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[27]) ? 1'b0 : force_valid[27];
assign force_wr_enable_splitted[30*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[72]) ? 1'b0 : force_valid[72];
assign force_wr_enable_splitted[30*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[82]) ? 1'b0 : force_valid[82];
assign force_wr_enable_splitted[30*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[102]) ? force_valid[102] : 1'b0;
assign force_wr_enable_splitted[30*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[131]) ? force_valid[131] : 1'b0;
assign force_wr_enable_splitted[30*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[136]) ? 1'b0 : force_valid[136];
assign force_wr_enable_splitted[30*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[191]) ? force_valid[191] : 1'b0;
assign force_wr_enable_splitted[30*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[209]) ? force_valid[209] : 1'b0;
assign force_wr_enable_splitted[30*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[210]) ? 1'b0 : force_valid[210];
assign force_wr_enable_splitted[30*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[245]) ? force_valid[245] : 1'b0;
assign force_wr_enable_splitted[30*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[297]) ? force_valid[297] : 1'b0;
assign force_wr_enable_splitted[30*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[305]) ? 1'b0 : force_valid[305];
assign force_wr_enable_splitted[30*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[316]) ? 1'b0 : force_valid[316];
assign force_wr_enable_splitted[30*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[330]) ? force_valid[330] : 1'b0;
assign force_wr_enable_splitted[31*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[6]) ? 1'b0 : force_valid[6];
assign force_wr_enable_splitted[31*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[61]) ? 1'b0 : force_valid[61];
assign force_wr_enable_splitted[31*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[79]) ? 1'b0 : force_valid[79];
assign force_wr_enable_splitted[31*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[109]) ? force_valid[109] : 1'b0;
assign force_wr_enable_splitted[31*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[115]) ? 1'b0 : force_valid[115];
assign force_wr_enable_splitted[31*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[138]) ? force_valid[138] : 1'b0;
assign force_wr_enable_splitted[31*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[170]) ? force_valid[170] : 1'b0;
assign force_wr_enable_splitted[31*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[216]) ? force_valid[216] : 1'b0;
assign force_wr_enable_splitted[31*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[217]) ? 1'b0 : force_valid[217];
assign force_wr_enable_splitted[31*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[224]) ? force_valid[224] : 1'b0;
assign force_wr_enable_splitted[31*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[284]) ? 1'b0 : force_valid[284];
assign force_wr_enable_splitted[31*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[304]) ? force_valid[304] : 1'b0;
assign force_wr_enable_splitted[31*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[309]) ? force_valid[309] : 1'b0;
assign force_wr_enable_splitted[31*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[323]) ? 1'b0 : force_valid[323];
assign force_wr_enable_splitted[32*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[116]) ? force_valid[116] : 1'b0;
assign force_wr_enable_splitted[32*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[153]) ? 1'b0 : force_valid[153];
assign force_wr_enable_splitted[32*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[198]) ? 1'b0 : force_valid[198];
assign force_wr_enable_splitted[32*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[208]) ? 1'b0 : force_valid[208];
assign force_wr_enable_splitted[32*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[224]) ? 1'b0 : force_valid[224];
assign force_wr_enable_splitted[32*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[251]) ? force_valid[251] : 1'b0;
assign force_wr_enable_splitted[32*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[257]) ? force_valid[257] : 1'b0;
assign force_wr_enable_splitted[32*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[262]) ? 1'b0 : force_valid[262];
assign force_wr_enable_splitted[32*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[317]) ? force_valid[317] : 1'b0;
assign force_wr_enable_splitted[32*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[344]) ? force_valid[344] : 1'b0;
assign force_wr_enable_splitted[32*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[358]) ? 1'b0 : force_valid[358];
assign force_wr_enable_splitted[32*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[371]) ? force_valid[371] : 1'b0;
assign force_wr_enable_splitted[32*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[423]) ? force_valid[423] : 1'b0;
assign force_wr_enable_splitted[32*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[431]) ? 1'b0 : force_valid[431];
assign force_wr_enable_splitted[33*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[123]) ? force_valid[123] : 1'b0;
assign force_wr_enable_splitted[33*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[160]) ? 1'b0 : force_valid[160];
assign force_wr_enable_splitted[33*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[205]) ? 1'b0 : force_valid[205];
assign force_wr_enable_splitted[33*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[215]) ? 1'b0 : force_valid[215];
assign force_wr_enable_splitted[33*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[230]) ? force_valid[230] : 1'b0;
assign force_wr_enable_splitted[33*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[231]) ? 1'b0 : force_valid[231];
assign force_wr_enable_splitted[33*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[264]) ? force_valid[264] : 1'b0;
assign force_wr_enable_splitted[33*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[269]) ? 1'b0 : force_valid[269];
assign force_wr_enable_splitted[33*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[324]) ? force_valid[324] : 1'b0;
assign force_wr_enable_splitted[33*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[337]) ? 1'b0 : force_valid[337];
assign force_wr_enable_splitted[33*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[351]) ? force_valid[351] : 1'b0;
assign force_wr_enable_splitted[33*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[378]) ? force_valid[378] : 1'b0;
assign force_wr_enable_splitted[33*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[430]) ? force_valid[430] : 1'b0;
assign force_wr_enable_splitted[33*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[438]) ? 1'b0 : force_valid[438];
assign force_wr_enable_splitted[34*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[130]) ? force_valid[130] : 1'b0;
assign force_wr_enable_splitted[34*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[167]) ? 1'b0 : force_valid[167];
assign force_wr_enable_splitted[34*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[212]) ? 1'b0 : force_valid[212];
assign force_wr_enable_splitted[34*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[222]) ? 1'b0 : force_valid[222];
assign force_wr_enable_splitted[34*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[237]) ? force_valid[237] : 1'b0;
assign force_wr_enable_splitted[34*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[238]) ? 1'b0 : force_valid[238];
assign force_wr_enable_splitted[34*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[271]) ? force_valid[271] : 1'b0;
assign force_wr_enable_splitted[34*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[276]) ? 1'b0 : force_valid[276];
assign force_wr_enable_splitted[34*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[331]) ? force_valid[331] : 1'b0;
assign force_wr_enable_splitted[34*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[344]) ? 1'b0 : force_valid[344];
assign force_wr_enable_splitted[34*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[358]) ? force_valid[358] : 1'b0;
assign force_wr_enable_splitted[34*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[385]) ? force_valid[385] : 1'b0;
assign force_wr_enable_splitted[34*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[437]) ? force_valid[437] : 1'b0;
assign force_wr_enable_splitted[34*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[445]) ? 1'b0 : force_valid[445];
assign force_wr_enable_splitted[35*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[137]) ? force_valid[137] : 1'b0;
assign force_wr_enable_splitted[35*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[146]) ? 1'b0 : force_valid[146];
assign force_wr_enable_splitted[35*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[201]) ? 1'b0 : force_valid[201];
assign force_wr_enable_splitted[35*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[219]) ? 1'b0 : force_valid[219];
assign force_wr_enable_splitted[35*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[244]) ? force_valid[244] : 1'b0;
assign force_wr_enable_splitted[35*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[245]) ? 1'b0 : force_valid[245];
assign force_wr_enable_splitted[35*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[255]) ? 1'b0 : force_valid[255];
assign force_wr_enable_splitted[35*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[278]) ? force_valid[278] : 1'b0;
assign force_wr_enable_splitted[35*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[310]) ? force_valid[310] : 1'b0;
assign force_wr_enable_splitted[35*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[337]) ? force_valid[337] : 1'b0;
assign force_wr_enable_splitted[35*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[351]) ? 1'b0 : force_valid[351];
assign force_wr_enable_splitted[35*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[364]) ? force_valid[364] : 1'b0;
assign force_wr_enable_splitted[35*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[424]) ? 1'b0 : force_valid[424];
assign force_wr_enable_splitted[35*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[444]) ? force_valid[444] : 1'b0;
assign force_wr_enable_splitted[36*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[114]) ? 1'b0 : force_valid[114];
assign force_wr_enable_splitted[36*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[124]) ? 1'b0 : force_valid[124];
assign force_wr_enable_splitted[36*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[144]) ? force_valid[144] : 1'b0;
assign force_wr_enable_splitted[36*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[181]) ? 1'b0 : force_valid[181];
assign force_wr_enable_splitted[36*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[233]) ? force_valid[233] : 1'b0;
assign force_wr_enable_splitted[36*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[252]) ? 1'b0 : force_valid[252];
assign force_wr_enable_splitted[36*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[279]) ? force_valid[279] : 1'b0;
assign force_wr_enable_splitted[36*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[285]) ? force_valid[285] : 1'b0;
assign force_wr_enable_splitted[36*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[290]) ? 1'b0 : force_valid[290];
assign force_wr_enable_splitted[36*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[339]) ? force_valid[339] : 1'b0;
assign force_wr_enable_splitted[36*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[347]) ? 1'b0 : force_valid[347];
assign force_wr_enable_splitted[36*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[372]) ? force_valid[372] : 1'b0;
assign force_wr_enable_splitted[36*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[386]) ? 1'b0 : force_valid[386];
assign force_wr_enable_splitted[36*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[399]) ? force_valid[399] : 1'b0;
assign force_wr_enable_splitted[37*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[121]) ? 1'b0 : force_valid[121];
assign force_wr_enable_splitted[37*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[131]) ? 1'b0 : force_valid[131];
assign force_wr_enable_splitted[37*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[151]) ? force_valid[151] : 1'b0;
assign force_wr_enable_splitted[37*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[188]) ? 1'b0 : force_valid[188];
assign force_wr_enable_splitted[37*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[240]) ? force_valid[240] : 1'b0;
assign force_wr_enable_splitted[37*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[258]) ? force_valid[258] : 1'b0;
assign force_wr_enable_splitted[37*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[259]) ? 1'b0 : force_valid[259];
assign force_wr_enable_splitted[37*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[292]) ? force_valid[292] : 1'b0;
assign force_wr_enable_splitted[37*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[297]) ? 1'b0 : force_valid[297];
assign force_wr_enable_splitted[37*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[346]) ? force_valid[346] : 1'b0;
assign force_wr_enable_splitted[37*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[354]) ? 1'b0 : force_valid[354];
assign force_wr_enable_splitted[37*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[365]) ? 1'b0 : force_valid[365];
assign force_wr_enable_splitted[37*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[379]) ? force_valid[379] : 1'b0;
assign force_wr_enable_splitted[37*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[406]) ? force_valid[406] : 1'b0;
assign force_wr_enable_splitted[38*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[128]) ? 1'b0 : force_valid[128];
assign force_wr_enable_splitted[38*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[138]) ? 1'b0 : force_valid[138];
assign force_wr_enable_splitted[38*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[158]) ? force_valid[158] : 1'b0;
assign force_wr_enable_splitted[38*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[195]) ? 1'b0 : force_valid[195];
assign force_wr_enable_splitted[38*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[247]) ? force_valid[247] : 1'b0;
assign force_wr_enable_splitted[38*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[265]) ? force_valid[265] : 1'b0;
assign force_wr_enable_splitted[38*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[266]) ? 1'b0 : force_valid[266];
assign force_wr_enable_splitted[38*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[299]) ? force_valid[299] : 1'b0;
assign force_wr_enable_splitted[38*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[304]) ? 1'b0 : force_valid[304];
assign force_wr_enable_splitted[38*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[353]) ? force_valid[353] : 1'b0;
assign force_wr_enable_splitted[38*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[361]) ? 1'b0 : force_valid[361];
assign force_wr_enable_splitted[38*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[372]) ? 1'b0 : force_valid[372];
assign force_wr_enable_splitted[38*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[386]) ? force_valid[386] : 1'b0;
assign force_wr_enable_splitted[38*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[413]) ? force_valid[413] : 1'b0;
assign force_wr_enable_splitted[39*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[117]) ? 1'b0 : force_valid[117];
assign force_wr_enable_splitted[39*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[135]) ? 1'b0 : force_valid[135];
assign force_wr_enable_splitted[39*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[165]) ? force_valid[165] : 1'b0;
assign force_wr_enable_splitted[39*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[174]) ? 1'b0 : force_valid[174];
assign force_wr_enable_splitted[39*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[226]) ? force_valid[226] : 1'b0;
assign force_wr_enable_splitted[39*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[272]) ? force_valid[272] : 1'b0;
assign force_wr_enable_splitted[39*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[273]) ? 1'b0 : force_valid[273];
assign force_wr_enable_splitted[39*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[283]) ? 1'b0 : force_valid[283];
assign force_wr_enable_splitted[39*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[306]) ? force_valid[306] : 1'b0;
assign force_wr_enable_splitted[39*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[340]) ? 1'b0 : force_valid[340];
assign force_wr_enable_splitted[39*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[360]) ? force_valid[360] : 1'b0;
assign force_wr_enable_splitted[39*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[365]) ? force_valid[365] : 1'b0;
assign force_wr_enable_splitted[39*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[379]) ? 1'b0 : force_valid[379];
assign force_wr_enable_splitted[39*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[392]) ? force_valid[392] : 1'b0;
assign force_wr_enable_splitted[40*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[142]) ? 1'b0 : force_valid[142];
assign force_wr_enable_splitted[40*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[152]) ? 1'b0 : force_valid[152];
assign force_wr_enable_splitted[40*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[172]) ? force_valid[172] : 1'b0;
assign force_wr_enable_splitted[40*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[209]) ? 1'b0 : force_valid[209];
assign force_wr_enable_splitted[40*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[261]) ? force_valid[261] : 1'b0;
assign force_wr_enable_splitted[40*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[280]) ? 1'b0 : force_valid[280];
assign force_wr_enable_splitted[40*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[307]) ? force_valid[307] : 1'b0;
assign force_wr_enable_splitted[40*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[313]) ? force_valid[313] : 1'b0;
assign force_wr_enable_splitted[40*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[318]) ? 1'b0 : force_valid[318];
assign force_wr_enable_splitted[40*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[367]) ? force_valid[367] : 1'b0;
assign force_wr_enable_splitted[40*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[375]) ? 1'b0 : force_valid[375];
assign force_wr_enable_splitted[40*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[400]) ? force_valid[400] : 1'b0;
assign force_wr_enable_splitted[40*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[414]) ? 1'b0 : force_valid[414];
assign force_wr_enable_splitted[40*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[427]) ? force_valid[427] : 1'b0;
assign force_wr_enable_splitted[41*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[149]) ? 1'b0 : force_valid[149];
assign force_wr_enable_splitted[41*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[159]) ? 1'b0 : force_valid[159];
assign force_wr_enable_splitted[41*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[179]) ? force_valid[179] : 1'b0;
assign force_wr_enable_splitted[41*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[216]) ? 1'b0 : force_valid[216];
assign force_wr_enable_splitted[41*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[268]) ? force_valid[268] : 1'b0;
assign force_wr_enable_splitted[41*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[286]) ? force_valid[286] : 1'b0;
assign force_wr_enable_splitted[41*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[287]) ? 1'b0 : force_valid[287];
assign force_wr_enable_splitted[41*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[320]) ? force_valid[320] : 1'b0;
assign force_wr_enable_splitted[41*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[325]) ? 1'b0 : force_valid[325];
assign force_wr_enable_splitted[41*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[374]) ? force_valid[374] : 1'b0;
assign force_wr_enable_splitted[41*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[382]) ? 1'b0 : force_valid[382];
assign force_wr_enable_splitted[41*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[393]) ? 1'b0 : force_valid[393];
assign force_wr_enable_splitted[41*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[407]) ? force_valid[407] : 1'b0;
assign force_wr_enable_splitted[41*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[434]) ? force_valid[434] : 1'b0;
assign force_wr_enable_splitted[42*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[156]) ? 1'b0 : force_valid[156];
assign force_wr_enable_splitted[42*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[166]) ? 1'b0 : force_valid[166];
assign force_wr_enable_splitted[42*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[186]) ? force_valid[186] : 1'b0;
assign force_wr_enable_splitted[42*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[223]) ? 1'b0 : force_valid[223];
assign force_wr_enable_splitted[42*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[275]) ? force_valid[275] : 1'b0;
assign force_wr_enable_splitted[42*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[293]) ? force_valid[293] : 1'b0;
assign force_wr_enable_splitted[42*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[294]) ? 1'b0 : force_valid[294];
assign force_wr_enable_splitted[42*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[327]) ? force_valid[327] : 1'b0;
assign force_wr_enable_splitted[42*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[332]) ? 1'b0 : force_valid[332];
assign force_wr_enable_splitted[42*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[381]) ? force_valid[381] : 1'b0;
assign force_wr_enable_splitted[42*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[389]) ? 1'b0 : force_valid[389];
assign force_wr_enable_splitted[42*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[400]) ? 1'b0 : force_valid[400];
assign force_wr_enable_splitted[42*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[414]) ? force_valid[414] : 1'b0;
assign force_wr_enable_splitted[42*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[441]) ? force_valid[441] : 1'b0;
assign force_wr_enable_splitted[43*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[145]) ? 1'b0 : force_valid[145];
assign force_wr_enable_splitted[43*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[163]) ? 1'b0 : force_valid[163];
assign force_wr_enable_splitted[43*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[193]) ? force_valid[193] : 1'b0;
assign force_wr_enable_splitted[43*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[202]) ? 1'b0 : force_valid[202];
assign force_wr_enable_splitted[43*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[254]) ? force_valid[254] : 1'b0;
assign force_wr_enable_splitted[43*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[300]) ? force_valid[300] : 1'b0;
assign force_wr_enable_splitted[43*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[301]) ? 1'b0 : force_valid[301];
assign force_wr_enable_splitted[43*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[311]) ? 1'b0 : force_valid[311];
assign force_wr_enable_splitted[43*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[334]) ? force_valid[334] : 1'b0;
assign force_wr_enable_splitted[43*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[368]) ? 1'b0 : force_valid[368];
assign force_wr_enable_splitted[43*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[388]) ? force_valid[388] : 1'b0;
assign force_wr_enable_splitted[43*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[393]) ? force_valid[393] : 1'b0;
assign force_wr_enable_splitted[43*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[407]) ? 1'b0 : force_valid[407];
assign force_wr_enable_splitted[43*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[420]) ? force_valid[420] : 1'b0;
assign force_wr_enable_splitted[44*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[125]) ? 1'b0 : force_valid[125];
assign force_wr_enable_splitted[44*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[170]) ? 1'b0 : force_valid[170];
assign force_wr_enable_splitted[44*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[180]) ? 1'b0 : force_valid[180];
assign force_wr_enable_splitted[44*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[200]) ? force_valid[200] : 1'b0;
assign force_wr_enable_splitted[44*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[229]) ? force_valid[229] : 1'b0;
assign force_wr_enable_splitted[44*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[234]) ? 1'b0 : force_valid[234];
assign force_wr_enable_splitted[44*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[289]) ? force_valid[289] : 1'b0;
assign force_wr_enable_splitted[44*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[308]) ? 1'b0 : force_valid[308];
assign force_wr_enable_splitted[44*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[335]) ? force_valid[335] : 1'b0;
assign force_wr_enable_splitted[44*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[343]) ? force_valid[343] : 1'b0;
assign force_wr_enable_splitted[44*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[395]) ? force_valid[395] : 1'b0;
assign force_wr_enable_splitted[44*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[403]) ? 1'b0 : force_valid[403];
assign force_wr_enable_splitted[44*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[428]) ? force_valid[428] : 1'b0;
assign force_wr_enable_splitted[44*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[442]) ? 1'b0 : force_valid[442];
assign force_wr_enable_splitted[45*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[132]) ? 1'b0 : force_valid[132];
assign force_wr_enable_splitted[45*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[177]) ? 1'b0 : force_valid[177];
assign force_wr_enable_splitted[45*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[187]) ? 1'b0 : force_valid[187];
assign force_wr_enable_splitted[45*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[207]) ? force_valid[207] : 1'b0;
assign force_wr_enable_splitted[45*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[236]) ? force_valid[236] : 1'b0;
assign force_wr_enable_splitted[45*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[241]) ? 1'b0 : force_valid[241];
assign force_wr_enable_splitted[45*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[296]) ? force_valid[296] : 1'b0;
assign force_wr_enable_splitted[45*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[314]) ? force_valid[314] : 1'b0;
assign force_wr_enable_splitted[45*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[315]) ? 1'b0 : force_valid[315];
assign force_wr_enable_splitted[45*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[350]) ? force_valid[350] : 1'b0;
assign force_wr_enable_splitted[45*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[402]) ? force_valid[402] : 1'b0;
assign force_wr_enable_splitted[45*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[410]) ? 1'b0 : force_valid[410];
assign force_wr_enable_splitted[45*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[421]) ? 1'b0 : force_valid[421];
assign force_wr_enable_splitted[45*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[435]) ? force_valid[435] : 1'b0;
assign force_wr_enable_splitted[46*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[139]) ? 1'b0 : force_valid[139];
assign force_wr_enable_splitted[46*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[184]) ? 1'b0 : force_valid[184];
assign force_wr_enable_splitted[46*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[194]) ? 1'b0 : force_valid[194];
assign force_wr_enable_splitted[46*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[214]) ? force_valid[214] : 1'b0;
assign force_wr_enable_splitted[46*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[243]) ? force_valid[243] : 1'b0;
assign force_wr_enable_splitted[46*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[248]) ? 1'b0 : force_valid[248];
assign force_wr_enable_splitted[46*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[303]) ? force_valid[303] : 1'b0;
assign force_wr_enable_splitted[46*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[321]) ? force_valid[321] : 1'b0;
assign force_wr_enable_splitted[46*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[322]) ? 1'b0 : force_valid[322];
assign force_wr_enable_splitted[46*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[357]) ? force_valid[357] : 1'b0;
assign force_wr_enable_splitted[46*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[409]) ? force_valid[409] : 1'b0;
assign force_wr_enable_splitted[46*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[417]) ? 1'b0 : force_valid[417];
assign force_wr_enable_splitted[46*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[428]) ? 1'b0 : force_valid[428];
assign force_wr_enable_splitted[46*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[442]) ? force_valid[442] : 1'b0;
assign force_wr_enable_splitted[47*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[118]) ? 1'b0 : force_valid[118];
assign force_wr_enable_splitted[47*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[173]) ? 1'b0 : force_valid[173];
assign force_wr_enable_splitted[47*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[191]) ? 1'b0 : force_valid[191];
assign force_wr_enable_splitted[47*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[221]) ? force_valid[221] : 1'b0;
assign force_wr_enable_splitted[47*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[227]) ? 1'b0 : force_valid[227];
assign force_wr_enable_splitted[47*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[250]) ? force_valid[250] : 1'b0;
assign force_wr_enable_splitted[47*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[282]) ? force_valid[282] : 1'b0;
assign force_wr_enable_splitted[47*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[328]) ? force_valid[328] : 1'b0;
assign force_wr_enable_splitted[47*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[329]) ? 1'b0 : force_valid[329];
assign force_wr_enable_splitted[47*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[336]) ? force_valid[336] : 1'b0;
assign force_wr_enable_splitted[47*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[396]) ? 1'b0 : force_valid[396];
assign force_wr_enable_splitted[47*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[416]) ? force_valid[416] : 1'b0;
assign force_wr_enable_splitted[47*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[421]) ? force_valid[421] : 1'b0;
assign force_wr_enable_splitted[47*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[435]) ? 1'b0 : force_valid[435];
assign force_wr_enable_splitted[48*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[8]) ? force_valid[8] : 1'b0;
assign force_wr_enable_splitted[48*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[22]) ? 1'b0 : force_valid[22];
assign force_wr_enable_splitted[48*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[35]) ? force_valid[35] : 1'b0;
assign force_wr_enable_splitted[48*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[87]) ? force_valid[87] : 1'b0;
assign force_wr_enable_splitted[48*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[95]) ? 1'b0 : force_valid[95];
assign force_wr_enable_splitted[48*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[228]) ? force_valid[228] : 1'b0;
assign force_wr_enable_splitted[48*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[265]) ? 1'b0 : force_valid[265];
assign force_wr_enable_splitted[48*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[310]) ? 1'b0 : force_valid[310];
assign force_wr_enable_splitted[48*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[320]) ? 1'b0 : force_valid[320];
assign force_wr_enable_splitted[48*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[336]) ? 1'b0 : force_valid[336];
assign force_wr_enable_splitted[48*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[363]) ? force_valid[363] : 1'b0;
assign force_wr_enable_splitted[48*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[369]) ? force_valid[369] : 1'b0;
assign force_wr_enable_splitted[48*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[374]) ? 1'b0 : force_valid[374];
assign force_wr_enable_splitted[48*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[429]) ? force_valid[429] : 1'b0;
assign force_wr_enable_splitted[49*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[1]) ? 1'b0 : force_valid[1];
assign force_wr_enable_splitted[49*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[15]) ? force_valid[15] : 1'b0;
assign force_wr_enable_splitted[49*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[42]) ? force_valid[42] : 1'b0;
assign force_wr_enable_splitted[49*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[94]) ? force_valid[94] : 1'b0;
assign force_wr_enable_splitted[49*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[102]) ? 1'b0 : force_valid[102];
assign force_wr_enable_splitted[49*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[235]) ? force_valid[235] : 1'b0;
assign force_wr_enable_splitted[49*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[272]) ? 1'b0 : force_valid[272];
assign force_wr_enable_splitted[49*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[317]) ? 1'b0 : force_valid[317];
assign force_wr_enable_splitted[49*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[327]) ? 1'b0 : force_valid[327];
assign force_wr_enable_splitted[49*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[342]) ? force_valid[342] : 1'b0;
assign force_wr_enable_splitted[49*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[343]) ? 1'b0 : force_valid[343];
assign force_wr_enable_splitted[49*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[376]) ? force_valid[376] : 1'b0;
assign force_wr_enable_splitted[49*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[381]) ? 1'b0 : force_valid[381];
assign force_wr_enable_splitted[49*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[436]) ? force_valid[436] : 1'b0;
assign force_wr_enable_splitted[50*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[8]) ? 1'b0 : force_valid[8];
assign force_wr_enable_splitted[50*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[22]) ? force_valid[22] : 1'b0;
assign force_wr_enable_splitted[50*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[49]) ? force_valid[49] : 1'b0;
assign force_wr_enable_splitted[50*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[101]) ? force_valid[101] : 1'b0;
assign force_wr_enable_splitted[50*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[109]) ? 1'b0 : force_valid[109];
assign force_wr_enable_splitted[50*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[242]) ? force_valid[242] : 1'b0;
assign force_wr_enable_splitted[50*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[279]) ? 1'b0 : force_valid[279];
assign force_wr_enable_splitted[50*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[324]) ? 1'b0 : force_valid[324];
assign force_wr_enable_splitted[50*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[334]) ? 1'b0 : force_valid[334];
assign force_wr_enable_splitted[50*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[349]) ? force_valid[349] : 1'b0;
assign force_wr_enable_splitted[50*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[350]) ? 1'b0 : force_valid[350];
assign force_wr_enable_splitted[50*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[383]) ? force_valid[383] : 1'b0;
assign force_wr_enable_splitted[50*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[388]) ? 1'b0 : force_valid[388];
assign force_wr_enable_splitted[50*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[443]) ? force_valid[443] : 1'b0;
assign force_wr_enable_splitted[51*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[1]) ? force_valid[1] : 1'b0;
assign force_wr_enable_splitted[51*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[15]) ? 1'b0 : force_valid[15];
assign force_wr_enable_splitted[51*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[28]) ? force_valid[28] : 1'b0;
assign force_wr_enable_splitted[51*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[88]) ? 1'b0 : force_valid[88];
assign force_wr_enable_splitted[51*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[108]) ? force_valid[108] : 1'b0;
assign force_wr_enable_splitted[51*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[249]) ? force_valid[249] : 1'b0;
assign force_wr_enable_splitted[51*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[258]) ? 1'b0 : force_valid[258];
assign force_wr_enable_splitted[51*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[313]) ? 1'b0 : force_valid[313];
assign force_wr_enable_splitted[51*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[331]) ? 1'b0 : force_valid[331];
assign force_wr_enable_splitted[51*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[356]) ? force_valid[356] : 1'b0;
assign force_wr_enable_splitted[51*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[357]) ? 1'b0 : force_valid[357];
assign force_wr_enable_splitted[51*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[367]) ? 1'b0 : force_valid[367];
assign force_wr_enable_splitted[51*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[390]) ? force_valid[390] : 1'b0;
assign force_wr_enable_splitted[51*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[422]) ? force_valid[422] : 1'b0;
assign force_wr_enable_splitted[52*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[3]) ? force_valid[3] : 1'b0;
assign force_wr_enable_splitted[52*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[11]) ? 1'b0 : force_valid[11];
assign force_wr_enable_splitted[52*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[36]) ? force_valid[36] : 1'b0;
assign force_wr_enable_splitted[52*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[50]) ? 1'b0 : force_valid[50];
assign force_wr_enable_splitted[52*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[63]) ? force_valid[63] : 1'b0;
assign force_wr_enable_splitted[52*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[226]) ? 1'b0 : force_valid[226];
assign force_wr_enable_splitted[52*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[236]) ? 1'b0 : force_valid[236];
assign force_wr_enable_splitted[52*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[256]) ? force_valid[256] : 1'b0;
assign force_wr_enable_splitted[52*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[293]) ? 1'b0 : force_valid[293];
assign force_wr_enable_splitted[52*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[345]) ? force_valid[345] : 1'b0;
assign force_wr_enable_splitted[52*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[364]) ? 1'b0 : force_valid[364];
assign force_wr_enable_splitted[52*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[391]) ? force_valid[391] : 1'b0;
assign force_wr_enable_splitted[52*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[397]) ? force_valid[397] : 1'b0;
assign force_wr_enable_splitted[52*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[402]) ? 1'b0 : force_valid[402];
assign force_wr_enable_splitted[53*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[10]) ? force_valid[10] : 1'b0;
assign force_wr_enable_splitted[53*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[18]) ? 1'b0 : force_valid[18];
assign force_wr_enable_splitted[53*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[29]) ? 1'b0 : force_valid[29];
assign force_wr_enable_splitted[53*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[43]) ? force_valid[43] : 1'b0;
assign force_wr_enable_splitted[53*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[70]) ? force_valid[70] : 1'b0;
assign force_wr_enable_splitted[53*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[233]) ? 1'b0 : force_valid[233];
assign force_wr_enable_splitted[53*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[243]) ? 1'b0 : force_valid[243];
assign force_wr_enable_splitted[53*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[263]) ? force_valid[263] : 1'b0;
assign force_wr_enable_splitted[53*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[300]) ? 1'b0 : force_valid[300];
assign force_wr_enable_splitted[53*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[352]) ? force_valid[352] : 1'b0;
assign force_wr_enable_splitted[53*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[370]) ? force_valid[370] : 1'b0;
assign force_wr_enable_splitted[53*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[371]) ? 1'b0 : force_valid[371];
assign force_wr_enable_splitted[53*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[404]) ? force_valid[404] : 1'b0;
assign force_wr_enable_splitted[53*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[409]) ? 1'b0 : force_valid[409];
assign force_wr_enable_splitted[54*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[17]) ? force_valid[17] : 1'b0;
assign force_wr_enable_splitted[54*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[25]) ? 1'b0 : force_valid[25];
assign force_wr_enable_splitted[54*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[36]) ? 1'b0 : force_valid[36];
assign force_wr_enable_splitted[54*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[50]) ? force_valid[50] : 1'b0;
assign force_wr_enable_splitted[54*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[77]) ? force_valid[77] : 1'b0;
assign force_wr_enable_splitted[54*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[240]) ? 1'b0 : force_valid[240];
assign force_wr_enable_splitted[54*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[250]) ? 1'b0 : force_valid[250];
assign force_wr_enable_splitted[54*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[270]) ? force_valid[270] : 1'b0;
assign force_wr_enable_splitted[54*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[307]) ? 1'b0 : force_valid[307];
assign force_wr_enable_splitted[54*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[359]) ? force_valid[359] : 1'b0;
assign force_wr_enable_splitted[54*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[377]) ? force_valid[377] : 1'b0;
assign force_wr_enable_splitted[54*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[378]) ? 1'b0 : force_valid[378];
assign force_wr_enable_splitted[54*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[411]) ? force_valid[411] : 1'b0;
assign force_wr_enable_splitted[54*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[416]) ? 1'b0 : force_valid[416];
assign force_wr_enable_splitted[55*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[4]) ? 1'b0 : force_valid[4];
assign force_wr_enable_splitted[55*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[24]) ? force_valid[24] : 1'b0;
assign force_wr_enable_splitted[55*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[29]) ? force_valid[29] : 1'b0;
assign force_wr_enable_splitted[55*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[43]) ? 1'b0 : force_valid[43];
assign force_wr_enable_splitted[55*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[56]) ? force_valid[56] : 1'b0;
assign force_wr_enable_splitted[55*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[229]) ? 1'b0 : force_valid[229];
assign force_wr_enable_splitted[55*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[247]) ? 1'b0 : force_valid[247];
assign force_wr_enable_splitted[55*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[277]) ? force_valid[277] : 1'b0;
assign force_wr_enable_splitted[55*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[286]) ? 1'b0 : force_valid[286];
assign force_wr_enable_splitted[55*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[338]) ? force_valid[338] : 1'b0;
assign force_wr_enable_splitted[55*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[384]) ? force_valid[384] : 1'b0;
assign force_wr_enable_splitted[55*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[385]) ? 1'b0 : force_valid[385];
assign force_wr_enable_splitted[55*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[395]) ? 1'b0 : force_valid[395];
assign force_wr_enable_splitted[55*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[418]) ? force_valid[418] : 1'b0;
assign force_wr_enable_splitted[56*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[31]) ? force_valid[31] : 1'b0;
assign force_wr_enable_splitted[56*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[39]) ? 1'b0 : force_valid[39];
assign force_wr_enable_splitted[56*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[64]) ? force_valid[64] : 1'b0;
assign force_wr_enable_splitted[56*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[78]) ? 1'b0 : force_valid[78];
assign force_wr_enable_splitted[56*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[91]) ? force_valid[91] : 1'b0;
assign force_wr_enable_splitted[56*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[254]) ? 1'b0 : force_valid[254];
assign force_wr_enable_splitted[56*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[264]) ? 1'b0 : force_valid[264];
assign force_wr_enable_splitted[56*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[284]) ? force_valid[284] : 1'b0;
assign force_wr_enable_splitted[56*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[321]) ? 1'b0 : force_valid[321];
assign force_wr_enable_splitted[56*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[373]) ? force_valid[373] : 1'b0;
assign force_wr_enable_splitted[56*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[392]) ? 1'b0 : force_valid[392];
assign force_wr_enable_splitted[56*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[419]) ? force_valid[419] : 1'b0;
assign force_wr_enable_splitted[56*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[425]) ? force_valid[425] : 1'b0;
assign force_wr_enable_splitted[56*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[430]) ? 1'b0 : force_valid[430];
assign force_wr_enable_splitted[57*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[38]) ? force_valid[38] : 1'b0;
assign force_wr_enable_splitted[57*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[46]) ? 1'b0 : force_valid[46];
assign force_wr_enable_splitted[57*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[57]) ? 1'b0 : force_valid[57];
assign force_wr_enable_splitted[57*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[71]) ? force_valid[71] : 1'b0;
assign force_wr_enable_splitted[57*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[98]) ? force_valid[98] : 1'b0;
assign force_wr_enable_splitted[57*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[261]) ? 1'b0 : force_valid[261];
assign force_wr_enable_splitted[57*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[271]) ? 1'b0 : force_valid[271];
assign force_wr_enable_splitted[57*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[291]) ? force_valid[291] : 1'b0;
assign force_wr_enable_splitted[57*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[328]) ? 1'b0 : force_valid[328];
assign force_wr_enable_splitted[57*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[380]) ? force_valid[380] : 1'b0;
assign force_wr_enable_splitted[57*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[398]) ? force_valid[398] : 1'b0;
assign force_wr_enable_splitted[57*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[399]) ? 1'b0 : force_valid[399];
assign force_wr_enable_splitted[57*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[432]) ? force_valid[432] : 1'b0;
assign force_wr_enable_splitted[57*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[437]) ? 1'b0 : force_valid[437];
assign force_wr_enable_splitted[58*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[45]) ? force_valid[45] : 1'b0;
assign force_wr_enable_splitted[58*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[53]) ? 1'b0 : force_valid[53];
assign force_wr_enable_splitted[58*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[64]) ? 1'b0 : force_valid[64];
assign force_wr_enable_splitted[58*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[78]) ? force_valid[78] : 1'b0;
assign force_wr_enable_splitted[58*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[105]) ? force_valid[105] : 1'b0;
assign force_wr_enable_splitted[58*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[268]) ? 1'b0 : force_valid[268];
assign force_wr_enable_splitted[58*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[278]) ? 1'b0 : force_valid[278];
assign force_wr_enable_splitted[58*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[298]) ? force_valid[298] : 1'b0;
assign force_wr_enable_splitted[58*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[335]) ? 1'b0 : force_valid[335];
assign force_wr_enable_splitted[58*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[387]) ? force_valid[387] : 1'b0;
assign force_wr_enable_splitted[58*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[405]) ? force_valid[405] : 1'b0;
assign force_wr_enable_splitted[58*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[406]) ? 1'b0 : force_valid[406];
assign force_wr_enable_splitted[58*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[439]) ? force_valid[439] : 1'b0;
assign force_wr_enable_splitted[58*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[444]) ? 1'b0 : force_valid[444];
assign force_wr_enable_splitted[59*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[32]) ? 1'b0 : force_valid[32];
assign force_wr_enable_splitted[59*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[52]) ? force_valid[52] : 1'b0;
assign force_wr_enable_splitted[59*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[57]) ? force_valid[57] : 1'b0;
assign force_wr_enable_splitted[59*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[71]) ? 1'b0 : force_valid[71];
assign force_wr_enable_splitted[59*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[84]) ? force_valid[84] : 1'b0;
assign force_wr_enable_splitted[59*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[257]) ? 1'b0 : force_valid[257];
assign force_wr_enable_splitted[59*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[275]) ? 1'b0 : force_valid[275];
assign force_wr_enable_splitted[59*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[305]) ? force_valid[305] : 1'b0;
assign force_wr_enable_splitted[59*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[314]) ? 1'b0 : force_valid[314];
assign force_wr_enable_splitted[59*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[366]) ? force_valid[366] : 1'b0;
assign force_wr_enable_splitted[59*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[412]) ? force_valid[412] : 1'b0;
assign force_wr_enable_splitted[59*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[413]) ? 1'b0 : force_valid[413];
assign force_wr_enable_splitted[59*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[423]) ? 1'b0 : force_valid[423];
assign force_wr_enable_splitted[59*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[446]) ? force_valid[446] : 1'b0;
assign force_wr_enable_splitted[60*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[7]) ? force_valid[7] : 1'b0;
assign force_wr_enable_splitted[60*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[59]) ? force_valid[59] : 1'b0;
assign force_wr_enable_splitted[60*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[67]) ? 1'b0 : force_valid[67];
assign force_wr_enable_splitted[60*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[92]) ? force_valid[92] : 1'b0;
assign force_wr_enable_splitted[60*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[106]) ? 1'b0 : force_valid[106];
assign force_wr_enable_splitted[60*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[237]) ? 1'b0 : force_valid[237];
assign force_wr_enable_splitted[60*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[282]) ? 1'b0 : force_valid[282];
assign force_wr_enable_splitted[60*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[292]) ? 1'b0 : force_valid[292];
assign force_wr_enable_splitted[60*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[312]) ? force_valid[312] : 1'b0;
assign force_wr_enable_splitted[60*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[341]) ? force_valid[341] : 1'b0;
assign force_wr_enable_splitted[60*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[346]) ? 1'b0 : force_valid[346];
assign force_wr_enable_splitted[60*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[401]) ? force_valid[401] : 1'b0;
assign force_wr_enable_splitted[60*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[420]) ? 1'b0 : force_valid[420];
assign force_wr_enable_splitted[60*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[447]) ? force_valid[447] : 1'b0;
assign force_wr_enable_splitted[61*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[14]) ? force_valid[14] : 1'b0;
assign force_wr_enable_splitted[61*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[66]) ? force_valid[66] : 1'b0;
assign force_wr_enable_splitted[61*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[74]) ? 1'b0 : force_valid[74];
assign force_wr_enable_splitted[61*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[85]) ? 1'b0 : force_valid[85];
assign force_wr_enable_splitted[61*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[99]) ? force_valid[99] : 1'b0;
assign force_wr_enable_splitted[61*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[244]) ? 1'b0 : force_valid[244];
assign force_wr_enable_splitted[61*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[289]) ? 1'b0 : force_valid[289];
assign force_wr_enable_splitted[61*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[299]) ? 1'b0 : force_valid[299];
assign force_wr_enable_splitted[61*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[319]) ? force_valid[319] : 1'b0;
assign force_wr_enable_splitted[61*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[348]) ? force_valid[348] : 1'b0;
assign force_wr_enable_splitted[61*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[353]) ? 1'b0 : force_valid[353];
assign force_wr_enable_splitted[61*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[408]) ? force_valid[408] : 1'b0;
assign force_wr_enable_splitted[61*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[426]) ? force_valid[426] : 1'b0;
assign force_wr_enable_splitted[61*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[427]) ? 1'b0 : force_valid[427];
assign force_wr_enable_splitted[62*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[21]) ? force_valid[21] : 1'b0;
assign force_wr_enable_splitted[62*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[73]) ? force_valid[73] : 1'b0;
assign force_wr_enable_splitted[62*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[81]) ? 1'b0 : force_valid[81];
assign force_wr_enable_splitted[62*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[92]) ? 1'b0 : force_valid[92];
assign force_wr_enable_splitted[62*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[106]) ? force_valid[106] : 1'b0;
assign force_wr_enable_splitted[62*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[251]) ? 1'b0 : force_valid[251];
assign force_wr_enable_splitted[62*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[296]) ? 1'b0 : force_valid[296];
assign force_wr_enable_splitted[62*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[306]) ? 1'b0 : force_valid[306];
assign force_wr_enable_splitted[62*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[326]) ? force_valid[326] : 1'b0;
assign force_wr_enable_splitted[62*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[355]) ? force_valid[355] : 1'b0;
assign force_wr_enable_splitted[62*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[360]) ? 1'b0 : force_valid[360];
assign force_wr_enable_splitted[62*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[415]) ? force_valid[415] : 1'b0;
assign force_wr_enable_splitted[62*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[433]) ? force_valid[433] : 1'b0;
assign force_wr_enable_splitted[62*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[434]) ? 1'b0 : force_valid[434];
assign force_wr_enable_splitted[63*(NUM_NEIGHBOR_CELLS+1)+0] = (force_dst[0]) ? force_valid[0] : 1'b0;
assign force_wr_enable_splitted[63*(NUM_NEIGHBOR_CELLS+1)+1] = (force_dst[60]) ? 1'b0 : force_valid[60];
assign force_wr_enable_splitted[63*(NUM_NEIGHBOR_CELLS+1)+2] = (force_dst[80]) ? force_valid[80] : 1'b0;
assign force_wr_enable_splitted[63*(NUM_NEIGHBOR_CELLS+1)+3] = (force_dst[85]) ? force_valid[85] : 1'b0;
assign force_wr_enable_splitted[63*(NUM_NEIGHBOR_CELLS+1)+4] = (force_dst[99]) ? 1'b0 : force_valid[99];
assign force_wr_enable_splitted[63*(NUM_NEIGHBOR_CELLS+1)+5] = (force_dst[230]) ? 1'b0 : force_valid[230];
assign force_wr_enable_splitted[63*(NUM_NEIGHBOR_CELLS+1)+6] = (force_dst[285]) ? 1'b0 : force_valid[285];
assign force_wr_enable_splitted[63*(NUM_NEIGHBOR_CELLS+1)+7] = (force_dst[303]) ? 1'b0 : force_valid[303];
assign force_wr_enable_splitted[63*(NUM_NEIGHBOR_CELLS+1)+8] = (force_dst[333]) ? force_valid[333] : 1'b0;
assign force_wr_enable_splitted[63*(NUM_NEIGHBOR_CELLS+1)+9] = (force_dst[339]) ? 1'b0 : force_valid[339];
assign force_wr_enable_splitted[63*(NUM_NEIGHBOR_CELLS+1)+10] = (force_dst[362]) ? force_valid[362] : 1'b0;
assign force_wr_enable_splitted[63*(NUM_NEIGHBOR_CELLS+1)+11] = (force_dst[394]) ? force_valid[394] : 1'b0;
assign force_wr_enable_splitted[63*(NUM_NEIGHBOR_CELLS+1)+12] = (force_dst[440]) ? force_valid[440] : 1'b0;
assign force_wr_enable_splitted[63*(NUM_NEIGHBOR_CELLS+1)+13] = (force_dst[441]) ? 1'b0 : force_valid[441];

endmodule