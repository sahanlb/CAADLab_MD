// INPUT_PLL.v

// Generated using ACDS version 18.0 219

`timescale 1 ps / 1 ps
module INPUT_PLL (
		output wire  locked,   //  locked.export
		output wire  outclk_0, // outclk0.clk
		input  wire  refclk,   //  refclk.clk
		input  wire  rst       //   reset.reset
	);

	INPUT_PLL_altera_iopll_180_ojuwjmy iopll_0 (
		.rst      (rst),      //   input,  width = 1,   reset.reset
		.refclk   (refclk),   //   input,  width = 1,  refclk.clk
		.locked   (locked),   //  output,  width = 1,  locked.export
		.outclk_0 (outclk_0)  //  output,  width = 1, outclk0.clk
	);

endmodule
