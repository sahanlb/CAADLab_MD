module all_position_caches
#(
	parameter NUM_CELLS = 64, 
	parameter DATA_WIDTH = 29, 
	parameter CELL_ID_WIDTH = 3,
	parameter NUM_PARTICLE_PER_CELL = 128, 
	parameter PARTICLE_ID_WIDTH = 7
)
(
	input clk,
	input rst,
	input Motion_Update_enable,
	input [PARTICLE_ID_WIDTH-1:0] MU_rd_addr,
	input [PARTICLE_ID_WIDTH-1:0] rd_addr,
	input [3*DATA_WIDTH-1:0] MU_wr_data,
	input [3*CELL_ID_WIDTH-1:0] MU_dst_cell,
	input MU_wr_data_valid,
	input MU_rden,
	
	output [NUM_CELLS*3*DATA_WIDTH-1:0] pos_data_out
);
	
	Pos_Cache_1_1_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(1)
	)
	cell_1_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[1*3*DATA_WIDTH-1:0*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_1_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(2)
	)
	cell_1_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[2*3*DATA_WIDTH-1:1*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_1_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(3)
	)
	cell_1_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[3*3*DATA_WIDTH-1:2*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_1_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(1),
		.CELL_Z(4)
	)
	cell_1_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[4*3*DATA_WIDTH-1:3*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_2_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(1)
	)
	cell_1_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[5*3*DATA_WIDTH-1:4*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(2)
	)
	cell_1_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[6*3*DATA_WIDTH-1:5*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_2_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(3)
	)
	cell_1_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[7*3*DATA_WIDTH-1:6*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_2_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(2),
		.CELL_Z(4)
	)
	cell_1_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[8*3*DATA_WIDTH-1:7*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_3_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(1)
	)
	cell_1_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[9*3*DATA_WIDTH-1:8*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_3_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(2)
	)
	cell_1_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[10*3*DATA_WIDTH-1:9*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_3_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(3)
	)
	cell_1_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[11*3*DATA_WIDTH-1:10*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_3_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(3),
		.CELL_Z(4)
	)
	cell_1_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[12*3*DATA_WIDTH-1:11*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_4_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(1)
	)
	cell_1_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[13*3*DATA_WIDTH-1:12*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_4_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(2)
	)
	cell_1_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[14*3*DATA_WIDTH-1:13*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_4_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(3)
	)
	cell_1_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[15*3*DATA_WIDTH-1:14*3*DATA_WIDTH])
	);
	
	Pos_Cache_1_4_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(1),
		.CELL_Y(4),
		.CELL_Z(4)
	)
	cell_1_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[16*3*DATA_WIDTH-1:15*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_1_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(1)
	)
	cell_2_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[17*3*DATA_WIDTH-1:16*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_1_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(2)
	)
	cell_2_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[18*3*DATA_WIDTH-1:17*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_1_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(3)
	)
	cell_2_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[19*3*DATA_WIDTH-1:18*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_1_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(1),
		.CELL_Z(4)
	)
	cell_2_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[20*3*DATA_WIDTH-1:19*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_2_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(1)
	)
	cell_2_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[21*3*DATA_WIDTH-1:20*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(2)
	)
	cell_2_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[22*3*DATA_WIDTH-1:21*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_2_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(3)
	)
	cell_2_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[23*3*DATA_WIDTH-1:22*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_2_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(2),
		.CELL_Z(4)
	)
	cell_2_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[24*3*DATA_WIDTH-1:23*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_3_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(1)
	)
	cell_2_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[25*3*DATA_WIDTH-1:24*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_3_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(2)
	)
	cell_2_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[26*3*DATA_WIDTH-1:25*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_3_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(3)
	)
	cell_2_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[27*3*DATA_WIDTH-1:26*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_3_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(3),
		.CELL_Z(4)
	)
	cell_2_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[28*3*DATA_WIDTH-1:27*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_4_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(1)
	)
	cell_2_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[29*3*DATA_WIDTH-1:28*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_4_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(2)
	)
	cell_2_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[30*3*DATA_WIDTH-1:29*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_4_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(3)
	)
	cell_2_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[31*3*DATA_WIDTH-1:30*3*DATA_WIDTH])
	);
	
	Pos_Cache_2_4_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(2),
		.CELL_Y(4),
		.CELL_Z(4)
	)
	cell_2_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[32*3*DATA_WIDTH-1:31*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_1_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(1)
	)
	cell_3_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[33*3*DATA_WIDTH-1:32*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_1_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(2)
	)
	cell_3_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[34*3*DATA_WIDTH-1:33*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_1_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(3)
	)
	cell_3_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[35*3*DATA_WIDTH-1:34*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_1_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(1),
		.CELL_Z(4)
	)
	cell_3_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[36*3*DATA_WIDTH-1:35*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_2_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(1)
	)
	cell_3_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[37*3*DATA_WIDTH-1:36*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(2)
	)
	cell_3_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[38*3*DATA_WIDTH-1:37*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_2_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(3)
	)
	cell_3_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[39*3*DATA_WIDTH-1:38*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_2_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(2),
		.CELL_Z(4)
	)
	cell_3_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[40*3*DATA_WIDTH-1:39*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_3_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(1)
	)
	cell_3_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[41*3*DATA_WIDTH-1:40*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_3_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(2)
	)
	cell_3_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[42*3*DATA_WIDTH-1:41*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_3_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(3)
	)
	cell_3_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[43*3*DATA_WIDTH-1:42*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_3_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(3),
		.CELL_Z(4)
	)
	cell_3_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[44*3*DATA_WIDTH-1:43*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_4_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(1)
	)
	cell_3_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[45*3*DATA_WIDTH-1:44*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_4_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(2)
	)
	cell_3_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[46*3*DATA_WIDTH-1:45*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_4_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(3)
	)
	cell_3_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[47*3*DATA_WIDTH-1:46*3*DATA_WIDTH])
	);
	
	Pos_Cache_3_4_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(3),
		.CELL_Y(4),
		.CELL_Z(4)
	)
	cell_3_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[48*3*DATA_WIDTH-1:47*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_1_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(1)
	)
	cell_4_1_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[49*3*DATA_WIDTH-1:48*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_1_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(2)
	)
	cell_4_1_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[50*3*DATA_WIDTH-1:49*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_1_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(3)
	)
	cell_4_1_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[51*3*DATA_WIDTH-1:50*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_1_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(1),
		.CELL_Z(4)
	)
	cell_4_1_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[52*3*DATA_WIDTH-1:51*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_2_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(1)
	)
	cell_4_2_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[53*3*DATA_WIDTH-1:52*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_2_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(2)
	)
	cell_4_2_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[54*3*DATA_WIDTH-1:53*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_2_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(3)
	)
	cell_4_2_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[55*3*DATA_WIDTH-1:54*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_2_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(2),
		.CELL_Z(4)
	)
	cell_4_2_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[56*3*DATA_WIDTH-1:55*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_3_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(1)
	)
	cell_4_3_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[57*3*DATA_WIDTH-1:56*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_3_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(2)
	)
	cell_4_3_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[58*3*DATA_WIDTH-1:57*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_3_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(3)
	)
	cell_4_3_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden :1'b1),
		.out_particle_info(pos_data_out[59*3*DATA_WIDTH-1:58*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_3_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(3),
		.CELL_Z(4)
	)
	cell_4_3_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[60*3*DATA_WIDTH-1:59*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_4_1
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(1)
	)
	cell_4_4_1
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[61*3*DATA_WIDTH-1:60*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_4_2
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(2)
	)
	cell_4_4_2
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[62*3*DATA_WIDTH-1:61*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_4_3
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(3)
	)
	cell_4_4_3
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[63*3*DATA_WIDTH-1:62*3*DATA_WIDTH])
	);
	
	Pos_Cache_4_4_4
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.PARTICLE_NUM(NUM_PARTICLE_PER_CELL),
		.ADDR_WIDTH(PARTICLE_ID_WIDTH),
		.CELL_ID_WIDTH(CELL_ID_WIDTH),
		.CELL_X(4),
		.CELL_Y(4),
		.CELL_Z(4)
	)
	cell_4_4_4
	(
		.clk(clk),
		.rst(rst),
		.motion_update_enable(Motion_Update_enable),				// Keep this signal as high during the motion update process
		.in_read_address(Motion_Update_enable ? MU_rd_addr : rd_addr),
		.in_data(MU_wr_data),
		.in_data_dst_cell(MU_dst_cell),				// The destination cell for the incoming data
		.in_data_valid(MU_wr_data_valid),						// Signify if the new incoming data is valid
		.in_rden(Motion_Update_enable ? MU_rden : 1'b1),
		.out_particle_info(pos_data_out[64*3*DATA_WIDTH-1:63*3*DATA_WIDTH])
	);
	
endmodule